module DCR(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [15:0] io_host_aw_bits_addr,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [31:0] io_host_w_bits_data,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [15:0] io_host_ar_bits_addr,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [31:0] io_host_r_bits_data,
  output        io_dcr_launch,
  input         io_dcr_finish,
  input         io_dcr_ecnt_0_valid,
  input  [31:0] io_dcr_ecnt_0_bits,
  output [31:0] io_dcr_ptrs_0,
  output [31:0] io_dcr_ptrs_1,
  output [31:0] io_dcr_ptrs_2,
  output [31:0] io_dcr_ptrs_3,
  output [31:0] io_dcr_ptrs_4,
  output [31:0] io_dcr_ptrs_5
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] waddr; // @[DCR.scala 88:22]
  reg [1:0] wstate; // @[DCR.scala 91:23]
  reg  rstate; // @[DCR.scala 95:23]
  reg [31:0] rdata; // @[DCR.scala 96:22]
  reg [31:0] reg_0; // @[DCR.scala 102:37]
  reg [31:0] reg_1; // @[DCR.scala 102:37]
  reg [31:0] reg_2; // @[DCR.scala 102:37]
  reg [31:0] reg_3; // @[DCR.scala 102:37]
  reg [31:0] reg_4; // @[DCR.scala 102:37]
  reg [31:0] reg_5; // @[DCR.scala 102:37]
  reg [31:0] reg_6; // @[DCR.scala 102:37]
  reg [31:0] reg_7; // @[DCR.scala 102:37]
  wire  _T = 2'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_1 = 2'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == wstate; // @[Conditional.scala 37:30]
  wire  _T_3 = io_host_aw_ready & io_host_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = ~rstate; // @[Conditional.scala 37:30]
  wire  _GEN_7 = io_host_ar_valid | rstate; // @[DCR.scala 138:30]
  wire  _T_11 = io_host_w_ready & io_host_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_12 = 16'h0 == waddr; // @[DCR.scala 156:44]
  wire  _T_13 = _T_11 & _T_12; // @[DCR.scala 156:31]
  wire  _T_15 = 16'h4 == waddr; // @[DCR.scala 163:51]
  wire  _T_16 = _T_11 & _T_15; // @[DCR.scala 163:33]
  wire  _T_18 = 16'h8 == waddr; // @[DCR.scala 169:45]
  wire  _T_19 = _T_11 & _T_18; // @[DCR.scala 169:27]
  wire  _T_21 = 16'hc == waddr; // @[DCR.scala 169:45]
  wire  _T_22 = _T_11 & _T_21; // @[DCR.scala 169:27]
  wire  _T_24 = 16'h10 == waddr; // @[DCR.scala 169:45]
  wire  _T_25 = _T_11 & _T_24; // @[DCR.scala 169:27]
  wire  _T_27 = 16'h14 == waddr; // @[DCR.scala 169:45]
  wire  _T_28 = _T_11 & _T_27; // @[DCR.scala 169:27]
  wire  _T_30 = 16'h18 == waddr; // @[DCR.scala 169:45]
  wire  _T_31 = _T_11 & _T_30; // @[DCR.scala 169:27]
  wire  _T_33 = 16'h1c == waddr; // @[DCR.scala 169:45]
  wire  _T_34 = _T_11 & _T_33; // @[DCR.scala 169:27]
  wire  _T_35 = io_host_ar_ready & io_host_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_36 = 16'h0 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_38 = 16'h4 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_40 = 16'h8 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_42 = 16'hc == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_44 = 16'h10 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_46 = 16'h14 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_48 = 16'h18 == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  wire  _T_50 = 16'h1c == io_host_ar_bits_addr; // @[Mux.scala 80:60]
  assign io_host_aw_ready = wstate == 2'h0; // @[DCR.scala 131:20]
  assign io_host_w_ready = wstate == 2'h1; // @[DCR.scala 132:19]
  assign io_host_b_valid = wstate == 2'h2; // @[DCR.scala 133:19]
  assign io_host_ar_ready = ~rstate; // @[DCR.scala 149:20]
  assign io_host_r_valid = rstate; // @[DCR.scala 150:19]
  assign io_host_r_bits_data = rdata; // @[DCR.scala 151:23]
  assign io_dcr_launch = reg_0[0]; // @[DCR.scala 178:17]
  assign io_dcr_ptrs_0 = reg_2; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_1 = reg_3; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_2 = reg_4; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_3 = reg_5; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_4 = reg_6; // @[DCR.scala 186:22]
  assign io_dcr_ptrs_5 = reg_7; // @[DCR.scala 186:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddr = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rstate = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  rdata = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_5 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_6 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_7 = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      waddr <= 16'hffff;
    end else if (_T_3) begin
      waddr <= io_host_aw_bits_addr;
    end
    if (reset) begin
      wstate <= 2'h0;
    end else if (_T) begin
      if (io_host_aw_valid) begin
        wstate <= 2'h1;
      end
    end else if (_T_1) begin
      if (io_host_w_valid) begin
        wstate <= 2'h2;
      end
    end else if (_T_2) begin
      if (io_host_b_ready) begin
        wstate <= 2'h0;
      end
    end
    if (reset) begin
      rstate <= 1'h0;
    end else if (_T_7) begin
      rstate <= _GEN_7;
    end else if (rstate) begin
      if (io_host_r_ready) begin
        rstate <= 1'h0;
      end
    end
    if (reset) begin
      rdata <= 32'h0;
    end else if (_T_35) begin
      if (_T_50) begin
        rdata <= reg_7;
      end else if (_T_48) begin
        rdata <= reg_6;
      end else if (_T_46) begin
        rdata <= reg_5;
      end else if (_T_44) begin
        rdata <= reg_4;
      end else if (_T_42) begin
        rdata <= reg_3;
      end else if (_T_40) begin
        rdata <= reg_2;
      end else if (_T_38) begin
        rdata <= reg_1;
      end else if (_T_36) begin
        rdata <= reg_0;
      end else begin
        rdata <= 32'h0;
      end
    end
    if (reset) begin
      reg_0 <= 32'h0;
    end else if (io_dcr_finish) begin
      reg_0 <= 32'h2;
    end else if (_T_13) begin
      reg_0 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_1 <= 32'h0;
    end else if (io_dcr_ecnt_0_valid) begin
      reg_1 <= io_dcr_ecnt_0_bits;
    end else if (_T_16) begin
      reg_1 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_2 <= 32'h0;
    end else if (_T_19) begin
      reg_2 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_3 <= 32'h0;
    end else if (_T_22) begin
      reg_3 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_4 <= 32'h0;
    end else if (_T_25) begin
      reg_4 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_5 <= 32'h0;
    end else if (_T_28) begin
      reg_5 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_6 <= 32'h0;
    end else if (_T_31) begin
      reg_6 <= io_host_w_bits_data;
    end
    if (reset) begin
      reg_7 <= 32'h0;
    end else if (_T_34) begin
      reg_7 <= io_host_w_bits_data;
    end
  end
endmodule
module Arbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
endmodule
module Arbiter_1(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [7:0]  io_in_1_bits_len,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [7:0]  io_in_2_bits_len,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [7:0]  io_in_3_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [7:0]  io_out_bits_len,
  output [1:0]  io_chosen
);
  wire [1:0] _GEN_0 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_1 = io_in_2_valid ? io_in_2_bits_len : io_in_3_bits_len; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_2 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_3 = io_in_1_valid ? 2'h1 : _GEN_0; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_4 = io_in_1_valid ? io_in_1_bits_len : _GEN_1; // @[Arbiter.scala 126:27]
  wire [31:0] _GEN_5 = io_in_1_valid ? io_in_1_bits_addr : _GEN_2; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  grant_2 = ~_T; // @[Arbiter.scala 31:78]
  wire  grant_3 = ~_T_1; // @[Arbiter.scala 31:78]
  wire  _T_6 = ~grant_3; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_2_ready = grant_2 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_3_ready = grant_3 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_6 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_5; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_len = io_in_0_valid ? 8'h7 : _GEN_4; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 2'h0 : _GEN_3; // @[Arbiter.scala 123:13 Arbiter.scala 127:17 Arbiter.scala 127:17 Arbiter.scala 127:17]
endmodule
module DME(
  input         clock,
  input         reset,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [7:0]  io_mem_aw_bits_len,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [7:0]  io_mem_ar_bits_len,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  output        io_dme_rd_0_cmd_ready,
  input         io_dme_rd_0_cmd_valid,
  input  [31:0] io_dme_rd_0_cmd_bits_addr,
  input         io_dme_rd_0_data_ready,
  output        io_dme_rd_0_data_valid,
  output [63:0] io_dme_rd_0_data_bits,
  output        io_dme_wr_0_cmd_ready,
  input         io_dme_wr_0_cmd_valid,
  input  [31:0] io_dme_wr_0_cmd_bits_addr,
  output        io_dme_wr_0_data_ready,
  input         io_dme_wr_0_data_valid,
  input  [63:0] io_dme_wr_0_data_bits,
  output        io_dme_wr_0_ack,
  output        io_dme_wr_1_cmd_ready,
  input         io_dme_wr_1_cmd_valid,
  input  [31:0] io_dme_wr_1_cmd_bits_addr,
  input  [7:0]  io_dme_wr_1_cmd_bits_len,
  output        io_dme_wr_1_data_ready,
  input         io_dme_wr_1_data_valid,
  input  [63:0] io_dme_wr_1_data_bits,
  output        io_dme_wr_1_ack,
  output        io_dme_wr_2_cmd_ready,
  input         io_dme_wr_2_cmd_valid,
  input  [31:0] io_dme_wr_2_cmd_bits_addr,
  input  [7:0]  io_dme_wr_2_cmd_bits_len,
  output        io_dme_wr_2_data_ready,
  input         io_dme_wr_2_data_valid,
  input  [63:0] io_dme_wr_2_data_bits,
  output        io_dme_wr_2_ack,
  output        io_dme_wr_3_cmd_ready,
  input         io_dme_wr_3_cmd_valid,
  input  [31:0] io_dme_wr_3_cmd_bits_addr,
  input  [7:0]  io_dme_wr_3_cmd_bits_len,
  output        io_dme_wr_3_data_ready,
  input         io_dme_wr_3_data_valid,
  input  [63:0] io_dme_wr_3_data_bits,
  output        io_dme_wr_3_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  rd_arb_io_in_0_ready; // @[DME.scala 130:22]
  wire  rd_arb_io_in_0_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_in_0_bits_addr; // @[DME.scala 130:22]
  wire  rd_arb_io_out_ready; // @[DME.scala 130:22]
  wire  rd_arb_io_out_valid; // @[DME.scala 130:22]
  wire [31:0] rd_arb_io_out_bits_addr; // @[DME.scala 130:22]
  wire  wr_arb_io_in_0_ready; // @[DME.scala 160:22]
  wire  wr_arb_io_in_0_valid; // @[DME.scala 160:22]
  wire [31:0] wr_arb_io_in_0_bits_addr; // @[DME.scala 160:22]
  wire  wr_arb_io_in_1_ready; // @[DME.scala 160:22]
  wire  wr_arb_io_in_1_valid; // @[DME.scala 160:22]
  wire [31:0] wr_arb_io_in_1_bits_addr; // @[DME.scala 160:22]
  wire [7:0] wr_arb_io_in_1_bits_len; // @[DME.scala 160:22]
  wire  wr_arb_io_in_2_ready; // @[DME.scala 160:22]
  wire  wr_arb_io_in_2_valid; // @[DME.scala 160:22]
  wire [31:0] wr_arb_io_in_2_bits_addr; // @[DME.scala 160:22]
  wire [7:0] wr_arb_io_in_2_bits_len; // @[DME.scala 160:22]
  wire  wr_arb_io_in_3_ready; // @[DME.scala 160:22]
  wire  wr_arb_io_in_3_valid; // @[DME.scala 160:22]
  wire [31:0] wr_arb_io_in_3_bits_addr; // @[DME.scala 160:22]
  wire [7:0] wr_arb_io_in_3_bits_len; // @[DME.scala 160:22]
  wire  wr_arb_io_out_ready; // @[DME.scala 160:22]
  wire  wr_arb_io_out_valid; // @[DME.scala 160:22]
  wire [31:0] wr_arb_io_out_bits_addr; // @[DME.scala 160:22]
  wire [7:0] wr_arb_io_out_bits_len; // @[DME.scala 160:22]
  wire [1:0] wr_arb_io_chosen; // @[DME.scala 160:22]
  wire  _T = rd_arb_io_out_ready & rd_arb_io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] rstate; // @[DME.scala 138:23]
  wire  _T_1 = 2'h0 == rstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == rstate; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == rstate; // @[Conditional.scala 37:30]
  wire  _T_4 = io_mem_r_ready & io_mem_r_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = _T_4 & io_mem_r_bits_last; // @[DME.scala 152:28]
  wire  _T_6 = wr_arb_io_out_ready & wr_arb_io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] wr_arb_chosen; // @[Reg.scala 15:16]
  reg [1:0] wstate; // @[DME.scala 168:23]
  reg [7:0] wr_cnt; // @[DME.scala 171:23]
  wire  _T_7 = wstate == 2'h0; // @[DME.scala 174:15]
  wire  _T_8 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 40:37]
  wire [7:0] _T_10 = wr_cnt + 8'h1; // @[DME.scala 177:22]
  wire  _T_11 = 2'h0 == wstate; // @[Conditional.scala 37:30]
  wire  _T_12 = 2'h1 == wstate; // @[Conditional.scala 37:30]
  wire  _T_13 = 2'h2 == wstate; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_23 = 2'h1 == wr_arb_chosen ? io_dme_wr_1_cmd_bits_len : 8'h7; // @[DME.scala 193:45]
  wire  _GEN_25 = 2'h1 == wr_arb_chosen ? io_dme_wr_1_data_valid : io_dme_wr_0_data_valid; // @[DME.scala 193:45]
  wire [63:0] _GEN_26 = 2'h1 == wr_arb_chosen ? io_dme_wr_1_data_bits : io_dme_wr_0_data_bits; // @[DME.scala 193:45]
  wire [7:0] _GEN_31 = 2'h2 == wr_arb_chosen ? io_dme_wr_2_cmd_bits_len : _GEN_23; // @[DME.scala 193:45]
  wire  _GEN_33 = 2'h2 == wr_arb_chosen ? io_dme_wr_2_data_valid : _GEN_25; // @[DME.scala 193:45]
  wire [63:0] _GEN_34 = 2'h2 == wr_arb_chosen ? io_dme_wr_2_data_bits : _GEN_26; // @[DME.scala 193:45]
  wire [7:0] _GEN_39 = 2'h3 == wr_arb_chosen ? io_dme_wr_3_cmd_bits_len : _GEN_31; // @[DME.scala 193:45]
  wire  _GEN_41 = 2'h3 == wr_arb_chosen ? io_dme_wr_3_data_valid : _GEN_33; // @[DME.scala 193:45]
  wire  _T_14 = _GEN_41 & io_mem_w_ready; // @[DME.scala 193:45]
  wire  _T_15 = wr_cnt == _GEN_39; // @[DME.scala 193:73]
  wire  _T_16 = _T_14 & _T_15; // @[DME.scala 193:63]
  wire  _T_17 = 2'h3 == wstate; // @[Conditional.scala 37:30]
  reg [7:0] rd_len; // @[Reg.scala 27:20]
  reg [31:0] rd_addr; // @[Reg.scala 27:20]
  reg [7:0] wr_len; // @[Reg.scala 27:20]
  reg [31:0] wr_addr; // @[Reg.scala 27:20]
  wire  _T_26 = wr_arb_chosen == 2'h0; // @[DME.scala 221:40]
  wire  _T_27 = io_mem_b_ready & io_mem_b_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = wstate == 2'h2; // @[DME.scala 222:67]
  wire  _T_31 = _T_26 & _T_30; // @[DME.scala 222:56]
  wire  _T_33 = wr_arb_chosen == 2'h1; // @[DME.scala 221:40]
  wire  _T_38 = _T_33 & _T_30; // @[DME.scala 222:56]
  wire  _T_40 = wr_arb_chosen == 2'h2; // @[DME.scala 221:40]
  wire  _T_45 = _T_40 & _T_30; // @[DME.scala 222:56]
  wire  _T_47 = wr_arb_chosen == 2'h3; // @[DME.scala 221:40]
  wire  _T_52 = _T_47 & _T_30; // @[DME.scala 222:56]
  wire  _T_60 = rstate == 2'h2; // @[DME.scala 240:28]
  Arbiter rd_arb ( // @[DME.scala 130:22]
    .io_in_0_ready(rd_arb_io_in_0_ready),
    .io_in_0_valid(rd_arb_io_in_0_valid),
    .io_in_0_bits_addr(rd_arb_io_in_0_bits_addr),
    .io_out_ready(rd_arb_io_out_ready),
    .io_out_valid(rd_arb_io_out_valid),
    .io_out_bits_addr(rd_arb_io_out_bits_addr)
  );
  Arbiter_1 wr_arb ( // @[DME.scala 160:22]
    .io_in_0_ready(wr_arb_io_in_0_ready),
    .io_in_0_valid(wr_arb_io_in_0_valid),
    .io_in_0_bits_addr(wr_arb_io_in_0_bits_addr),
    .io_in_1_ready(wr_arb_io_in_1_ready),
    .io_in_1_valid(wr_arb_io_in_1_valid),
    .io_in_1_bits_addr(wr_arb_io_in_1_bits_addr),
    .io_in_1_bits_len(wr_arb_io_in_1_bits_len),
    .io_in_2_ready(wr_arb_io_in_2_ready),
    .io_in_2_valid(wr_arb_io_in_2_valid),
    .io_in_2_bits_addr(wr_arb_io_in_2_bits_addr),
    .io_in_2_bits_len(wr_arb_io_in_2_bits_len),
    .io_in_3_ready(wr_arb_io_in_3_ready),
    .io_in_3_valid(wr_arb_io_in_3_valid),
    .io_in_3_bits_addr(wr_arb_io_in_3_bits_addr),
    .io_in_3_bits_len(wr_arb_io_in_3_bits_len),
    .io_out_ready(wr_arb_io_out_ready),
    .io_out_valid(wr_arb_io_out_valid),
    .io_out_bits_addr(wr_arb_io_out_bits_addr),
    .io_out_bits_len(wr_arb_io_out_bits_len),
    .io_chosen(wr_arb_io_chosen)
  );
  assign io_mem_aw_valid = wstate == 2'h1; // @[DME.scala 226:19]
  assign io_mem_aw_bits_addr = wr_addr; // @[DME.scala 227:23]
  assign io_mem_aw_bits_len = wr_len; // @[DME.scala 228:22]
  assign io_mem_w_valid = _T_30 & _GEN_41; // @[DME.scala 230:18]
  assign io_mem_w_bits_data = 2'h3 == wr_arb_chosen ? io_dme_wr_3_data_bits : _GEN_34; // @[DME.scala 231:22]
  assign io_mem_w_bits_last = wr_cnt == _GEN_39; // @[DME.scala 232:22]
  assign io_mem_b_ready = wstate == 2'h3; // @[DME.scala 234:18]
  assign io_mem_ar_valid = rstate == 2'h1; // @[DME.scala 236:19]
  assign io_mem_ar_bits_addr = rd_addr; // @[DME.scala 237:23]
  assign io_mem_ar_bits_len = rd_len; // @[DME.scala 238:22]
  assign io_mem_r_ready = _T_60 & io_dme_rd_0_data_ready; // @[DME.scala 240:18]
  assign io_dme_rd_0_cmd_ready = rd_arb_io_in_0_ready; // @[DME.scala 134:21]
  assign io_dme_rd_0_data_valid = io_mem_r_valid; // @[DME.scala 215:29]
  assign io_dme_rd_0_data_bits = io_mem_r_bits_data; // @[DME.scala 216:28]
  assign io_dme_wr_0_cmd_ready = wr_arb_io_in_0_ready; // @[DME.scala 164:21]
  assign io_dme_wr_0_data_ready = _T_31 & io_mem_w_ready; // @[DME.scala 222:29]
  assign io_dme_wr_0_ack = _T_26 & _T_27; // @[DME.scala 221:22]
  assign io_dme_wr_1_cmd_ready = wr_arb_io_in_1_ready; // @[DME.scala 164:21]
  assign io_dme_wr_1_data_ready = _T_38 & io_mem_w_ready; // @[DME.scala 222:29]
  assign io_dme_wr_1_ack = _T_33 & _T_27; // @[DME.scala 221:22]
  assign io_dme_wr_2_cmd_ready = wr_arb_io_in_2_ready; // @[DME.scala 164:21]
  assign io_dme_wr_2_data_ready = _T_45 & io_mem_w_ready; // @[DME.scala 222:29]
  assign io_dme_wr_2_ack = _T_40 & _T_27; // @[DME.scala 221:22]
  assign io_dme_wr_3_cmd_ready = wr_arb_io_in_3_ready; // @[DME.scala 164:21]
  assign io_dme_wr_3_data_ready = _T_52 & io_mem_w_ready; // @[DME.scala 222:29]
  assign io_dme_wr_3_ack = _T_47 & _T_27; // @[DME.scala 221:22]
  assign rd_arb_io_in_0_valid = io_dme_rd_0_cmd_valid; // @[DME.scala 134:21]
  assign rd_arb_io_in_0_bits_addr = io_dme_rd_0_cmd_bits_addr; // @[DME.scala 134:21]
  assign rd_arb_io_out_ready = rstate == 2'h0; // @[DME.scala 210:23]
  assign wr_arb_io_in_0_valid = io_dme_wr_0_cmd_valid; // @[DME.scala 164:21]
  assign wr_arb_io_in_0_bits_addr = io_dme_wr_0_cmd_bits_addr; // @[DME.scala 164:21]
  assign wr_arb_io_in_1_valid = io_dme_wr_1_cmd_valid; // @[DME.scala 164:21]
  assign wr_arb_io_in_1_bits_addr = io_dme_wr_1_cmd_bits_addr; // @[DME.scala 164:21]
  assign wr_arb_io_in_1_bits_len = io_dme_wr_1_cmd_bits_len; // @[DME.scala 164:21]
  assign wr_arb_io_in_2_valid = io_dme_wr_2_cmd_valid; // @[DME.scala 164:21]
  assign wr_arb_io_in_2_bits_addr = io_dme_wr_2_cmd_bits_addr; // @[DME.scala 164:21]
  assign wr_arb_io_in_2_bits_len = io_dme_wr_2_cmd_bits_len; // @[DME.scala 164:21]
  assign wr_arb_io_in_3_valid = io_dme_wr_3_cmd_valid; // @[DME.scala 164:21]
  assign wr_arb_io_in_3_bits_addr = io_dme_wr_3_cmd_bits_addr; // @[DME.scala 164:21]
  assign wr_arb_io_in_3_bits_len = io_dme_wr_3_cmd_bits_len; // @[DME.scala 164:21]
  assign wr_arb_io_out_ready = wstate == 2'h0; // @[DME.scala 211:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rstate = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  wr_arb_chosen = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  wstate = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  wr_cnt = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  rd_len = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  rd_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  wr_len = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  wr_addr = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      rstate <= 2'h0;
    end else if (_T_1) begin
      if (rd_arb_io_out_valid) begin
        rstate <= 2'h1;
      end
    end else if (_T_2) begin
      if (io_mem_ar_ready) begin
        rstate <= 2'h2;
      end
    end else if (_T_3) begin
      if (_T_5) begin
        rstate <= 2'h0;
      end
    end
    if (_T_6) begin
      wr_arb_chosen <= wr_arb_io_chosen;
    end
    if (reset) begin
      wstate <= 2'h0;
    end else if (_T_11) begin
      if (wr_arb_io_out_valid) begin
        wstate <= 2'h1;
      end
    end else if (_T_12) begin
      if (io_mem_aw_ready) begin
        wstate <= 2'h2;
      end
    end else if (_T_13) begin
      if (_T_16) begin
        wstate <= 2'h3;
      end
    end else if (_T_17) begin
      if (io_mem_b_valid) begin
        wstate <= 2'h0;
      end
    end
    if (reset) begin
      wr_cnt <= 8'h0;
    end else if (_T_7) begin
      wr_cnt <= 8'h0;
    end else if (_T_8) begin
      wr_cnt <= _T_10;
    end
    if (reset) begin
      rd_len <= 8'h0;
    end else if (_T) begin
      rd_len <= 8'h7;
    end
    if (reset) begin
      rd_addr <= 32'h0;
    end else if (_T) begin
      rd_addr <= rd_arb_io_out_bits_addr;
    end
    if (reset) begin
      wr_len <= 8'h0;
    end else if (_T_6) begin
      wr_len <= wr_arb_io_out_bits_len;
    end
    if (reset) begin
      wr_addr <= 32'h0;
    end else if (_T_6) begin
      wr_addr <= wr_arb_io_out_bits_addr;
    end
  end
endmodule
module DMECache(
  input         clock,
  input         reset,
  input         io_cpu_flush,
  output        io_cpu_flush_done,
  output        io_cpu_req_ready,
  input         io_cpu_req_valid,
  input  [63:0] io_cpu_req_bits_addr,
  input  [63:0] io_cpu_req_bits_data,
  input  [7:0]  io_cpu_req_bits_mask,
  input  [7:0]  io_cpu_req_bits_tag,
  output        io_cpu_resp_valid,
  output [63:0] io_cpu_resp_bits_data,
  output [7:0]  io_cpu_resp_bits_tag,
  input         io_mem_rd_cmd_ready,
  output        io_mem_rd_cmd_valid,
  output [31:0] io_mem_rd_cmd_bits_addr,
  output        io_mem_rd_data_ready,
  input         io_mem_rd_data_valid,
  input  [63:0] io_mem_rd_data_bits,
  input         io_mem_wr_cmd_ready,
  output        io_mem_wr_cmd_valid,
  output [31:0] io_mem_wr_cmd_bits_addr,
  input         io_mem_wr_data_ready,
  output        io_mem_wr_data_valid,
  output [63:0] io_mem_wr_data_bits,
  input         io_mem_wr_ack
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_257;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [255:0] _RAND_264;
  reg [255:0] _RAND_265;
  reg [63:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [63:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [63:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [511:0] _RAND_276;
  reg [63:0] _RAND_277;
  reg [63:0] _RAND_278;
  reg [63:0] _RAND_279;
  reg [63:0] _RAND_280;
  reg [63:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [63:0] _RAND_283;
  reg [63:0] _RAND_284;
`endif // RANDOMIZE_REG_INIT
  reg [49:0] metaMem_tag [0:255]; // @[AXICache.scala 720:28]
  wire [49:0] metaMem_tag_rmeta_data; // @[AXICache.scala 720:28]
  wire [7:0] metaMem_tag_rmeta_addr; // @[AXICache.scala 720:28]
  wire [49:0] metaMem_tag__T_431_data; // @[AXICache.scala 720:28]
  wire [7:0] metaMem_tag__T_431_addr; // @[AXICache.scala 720:28]
  wire [49:0] metaMem_tag__T_262_data; // @[AXICache.scala 720:28]
  wire [7:0] metaMem_tag__T_262_addr; // @[AXICache.scala 720:28]
  wire  metaMem_tag__T_262_mask; // @[AXICache.scala 720:28]
  wire  metaMem_tag__T_262_en; // @[AXICache.scala 720:28]
  reg  metaMem_tag_rmeta_en_pipe_0;
  reg [7:0] metaMem_tag_rmeta_addr_pipe_0;
  reg  metaMem_tag__T_431_en_pipe_0;
  reg [7:0] metaMem_tag__T_431_addr_pipe_0;
  reg [7:0] dataMem_0_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_0__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_0__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_0__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_0__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_0__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_0__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_0__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_0__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_0__T_14_addr_pipe_0;
  reg  dataMem_0_0__T_112_en_pipe_0;
  reg [7:0] dataMem_0_0__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_1__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_1__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_1__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_1__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_1__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_1__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_1__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_1__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_1__T_14_addr_pipe_0;
  reg  dataMem_0_1__T_112_en_pipe_0;
  reg [7:0] dataMem_0_1__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_2__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_2__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_2__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_2__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_2__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_2__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_2__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_2__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_2__T_14_addr_pipe_0;
  reg  dataMem_0_2__T_112_en_pipe_0;
  reg [7:0] dataMem_0_2__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_3__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_3__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_3__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_3__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_3__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_3__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_3__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_3__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_3__T_14_addr_pipe_0;
  reg  dataMem_0_3__T_112_en_pipe_0;
  reg [7:0] dataMem_0_3__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_4__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_4__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_4__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_4__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_4__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_4__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_4__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_4__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_4__T_14_addr_pipe_0;
  reg  dataMem_0_4__T_112_en_pipe_0;
  reg [7:0] dataMem_0_4__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_5__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_5__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_5__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_5__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_5__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_5__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_5__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_5__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_5__T_14_addr_pipe_0;
  reg  dataMem_0_5__T_112_en_pipe_0;
  reg [7:0] dataMem_0_5__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_6__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_6__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_6__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_6__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_6__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_6__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_6__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_6__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_6__T_14_addr_pipe_0;
  reg  dataMem_0_6__T_112_en_pipe_0;
  reg [7:0] dataMem_0_6__T_112_addr_pipe_0;
  reg [7:0] dataMem_0_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_7__T_14_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_7__T_14_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_7__T_112_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_7__T_112_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_7__T_281_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_0_7__T_281_addr; // @[AXICache.scala 721:45]
  wire  dataMem_0_7__T_281_mask; // @[AXICache.scala 721:45]
  wire  dataMem_0_7__T_281_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_0_7__T_14_addr_pipe_0;
  reg  dataMem_0_7__T_112_en_pipe_0;
  reg [7:0] dataMem_0_7__T_112_addr_pipe_0;
  reg [7:0] dataMem_1_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_0__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_0__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_0__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_0__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_0__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_0__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_0__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_0__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_0__T_24_addr_pipe_0;
  reg  dataMem_1_0__T_123_en_pipe_0;
  reg [7:0] dataMem_1_0__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_1__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_1__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_1__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_1__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_1__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_1__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_1__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_1__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_1__T_24_addr_pipe_0;
  reg  dataMem_1_1__T_123_en_pipe_0;
  reg [7:0] dataMem_1_1__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_2__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_2__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_2__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_2__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_2__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_2__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_2__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_2__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_2__T_24_addr_pipe_0;
  reg  dataMem_1_2__T_123_en_pipe_0;
  reg [7:0] dataMem_1_2__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_3__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_3__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_3__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_3__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_3__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_3__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_3__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_3__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_3__T_24_addr_pipe_0;
  reg  dataMem_1_3__T_123_en_pipe_0;
  reg [7:0] dataMem_1_3__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_4__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_4__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_4__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_4__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_4__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_4__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_4__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_4__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_4__T_24_addr_pipe_0;
  reg  dataMem_1_4__T_123_en_pipe_0;
  reg [7:0] dataMem_1_4__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_5__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_5__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_5__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_5__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_5__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_5__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_5__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_5__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_5__T_24_addr_pipe_0;
  reg  dataMem_1_5__T_123_en_pipe_0;
  reg [7:0] dataMem_1_5__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_6__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_6__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_6__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_6__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_6__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_6__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_6__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_6__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_6__T_24_addr_pipe_0;
  reg  dataMem_1_6__T_123_en_pipe_0;
  reg [7:0] dataMem_1_6__T_123_addr_pipe_0;
  reg [7:0] dataMem_1_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_7__T_24_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_7__T_24_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_7__T_123_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_7__T_123_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_7__T_300_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_1_7__T_300_addr; // @[AXICache.scala 721:45]
  wire  dataMem_1_7__T_300_mask; // @[AXICache.scala 721:45]
  wire  dataMem_1_7__T_300_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_1_7__T_24_addr_pipe_0;
  reg  dataMem_1_7__T_123_en_pipe_0;
  reg [7:0] dataMem_1_7__T_123_addr_pipe_0;
  reg [7:0] dataMem_2_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_0__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_0__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_0__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_0__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_0__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_0__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_0__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_0__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_0__T_34_addr_pipe_0;
  reg  dataMem_2_0__T_134_en_pipe_0;
  reg [7:0] dataMem_2_0__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_1__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_1__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_1__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_1__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_1__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_1__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_1__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_1__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_1__T_34_addr_pipe_0;
  reg  dataMem_2_1__T_134_en_pipe_0;
  reg [7:0] dataMem_2_1__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_2__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_2__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_2__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_2__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_2__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_2__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_2__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_2__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_2__T_34_addr_pipe_0;
  reg  dataMem_2_2__T_134_en_pipe_0;
  reg [7:0] dataMem_2_2__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_3__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_3__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_3__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_3__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_3__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_3__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_3__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_3__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_3__T_34_addr_pipe_0;
  reg  dataMem_2_3__T_134_en_pipe_0;
  reg [7:0] dataMem_2_3__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_4__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_4__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_4__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_4__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_4__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_4__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_4__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_4__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_4__T_34_addr_pipe_0;
  reg  dataMem_2_4__T_134_en_pipe_0;
  reg [7:0] dataMem_2_4__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_5__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_5__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_5__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_5__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_5__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_5__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_5__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_5__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_5__T_34_addr_pipe_0;
  reg  dataMem_2_5__T_134_en_pipe_0;
  reg [7:0] dataMem_2_5__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_6__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_6__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_6__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_6__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_6__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_6__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_6__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_6__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_6__T_34_addr_pipe_0;
  reg  dataMem_2_6__T_134_en_pipe_0;
  reg [7:0] dataMem_2_6__T_134_addr_pipe_0;
  reg [7:0] dataMem_2_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_7__T_34_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_7__T_34_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_7__T_134_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_7__T_134_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_7__T_319_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_2_7__T_319_addr; // @[AXICache.scala 721:45]
  wire  dataMem_2_7__T_319_mask; // @[AXICache.scala 721:45]
  wire  dataMem_2_7__T_319_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_2_7__T_34_addr_pipe_0;
  reg  dataMem_2_7__T_134_en_pipe_0;
  reg [7:0] dataMem_2_7__T_134_addr_pipe_0;
  reg [7:0] dataMem_3_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_0__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_0__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_0__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_0__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_0__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_0__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_0__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_0__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_0__T_44_addr_pipe_0;
  reg  dataMem_3_0__T_145_en_pipe_0;
  reg [7:0] dataMem_3_0__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_1__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_1__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_1__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_1__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_1__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_1__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_1__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_1__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_1__T_44_addr_pipe_0;
  reg  dataMem_3_1__T_145_en_pipe_0;
  reg [7:0] dataMem_3_1__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_2__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_2__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_2__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_2__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_2__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_2__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_2__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_2__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_2__T_44_addr_pipe_0;
  reg  dataMem_3_2__T_145_en_pipe_0;
  reg [7:0] dataMem_3_2__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_3__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_3__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_3__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_3__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_3__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_3__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_3__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_3__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_3__T_44_addr_pipe_0;
  reg  dataMem_3_3__T_145_en_pipe_0;
  reg [7:0] dataMem_3_3__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_4__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_4__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_4__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_4__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_4__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_4__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_4__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_4__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_4__T_44_addr_pipe_0;
  reg  dataMem_3_4__T_145_en_pipe_0;
  reg [7:0] dataMem_3_4__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_5__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_5__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_5__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_5__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_5__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_5__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_5__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_5__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_5__T_44_addr_pipe_0;
  reg  dataMem_3_5__T_145_en_pipe_0;
  reg [7:0] dataMem_3_5__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_6__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_6__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_6__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_6__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_6__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_6__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_6__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_6__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_6__T_44_addr_pipe_0;
  reg  dataMem_3_6__T_145_en_pipe_0;
  reg [7:0] dataMem_3_6__T_145_addr_pipe_0;
  reg [7:0] dataMem_3_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_7__T_44_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_7__T_44_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_7__T_145_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_7__T_145_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_7__T_338_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_3_7__T_338_addr; // @[AXICache.scala 721:45]
  wire  dataMem_3_7__T_338_mask; // @[AXICache.scala 721:45]
  wire  dataMem_3_7__T_338_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_3_7__T_44_addr_pipe_0;
  reg  dataMem_3_7__T_145_en_pipe_0;
  reg [7:0] dataMem_3_7__T_145_addr_pipe_0;
  reg [7:0] dataMem_4_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_0__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_0__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_0__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_0__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_0__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_0__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_0__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_0__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_0__T_54_addr_pipe_0;
  reg  dataMem_4_0__T_156_en_pipe_0;
  reg [7:0] dataMem_4_0__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_1__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_1__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_1__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_1__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_1__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_1__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_1__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_1__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_1__T_54_addr_pipe_0;
  reg  dataMem_4_1__T_156_en_pipe_0;
  reg [7:0] dataMem_4_1__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_2__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_2__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_2__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_2__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_2__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_2__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_2__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_2__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_2__T_54_addr_pipe_0;
  reg  dataMem_4_2__T_156_en_pipe_0;
  reg [7:0] dataMem_4_2__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_3__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_3__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_3__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_3__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_3__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_3__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_3__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_3__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_3__T_54_addr_pipe_0;
  reg  dataMem_4_3__T_156_en_pipe_0;
  reg [7:0] dataMem_4_3__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_4__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_4__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_4__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_4__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_4__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_4__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_4__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_4__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_4__T_54_addr_pipe_0;
  reg  dataMem_4_4__T_156_en_pipe_0;
  reg [7:0] dataMem_4_4__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_5__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_5__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_5__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_5__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_5__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_5__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_5__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_5__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_5__T_54_addr_pipe_0;
  reg  dataMem_4_5__T_156_en_pipe_0;
  reg [7:0] dataMem_4_5__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_6__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_6__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_6__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_6__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_6__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_6__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_6__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_6__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_6__T_54_addr_pipe_0;
  reg  dataMem_4_6__T_156_en_pipe_0;
  reg [7:0] dataMem_4_6__T_156_addr_pipe_0;
  reg [7:0] dataMem_4_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_7__T_54_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_7__T_54_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_7__T_156_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_7__T_156_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_7__T_357_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_4_7__T_357_addr; // @[AXICache.scala 721:45]
  wire  dataMem_4_7__T_357_mask; // @[AXICache.scala 721:45]
  wire  dataMem_4_7__T_357_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_4_7__T_54_addr_pipe_0;
  reg  dataMem_4_7__T_156_en_pipe_0;
  reg [7:0] dataMem_4_7__T_156_addr_pipe_0;
  reg [7:0] dataMem_5_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_0__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_0__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_0__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_0__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_0__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_0__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_0__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_0__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_0__T_64_addr_pipe_0;
  reg  dataMem_5_0__T_167_en_pipe_0;
  reg [7:0] dataMem_5_0__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_1__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_1__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_1__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_1__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_1__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_1__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_1__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_1__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_1__T_64_addr_pipe_0;
  reg  dataMem_5_1__T_167_en_pipe_0;
  reg [7:0] dataMem_5_1__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_2__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_2__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_2__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_2__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_2__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_2__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_2__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_2__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_2__T_64_addr_pipe_0;
  reg  dataMem_5_2__T_167_en_pipe_0;
  reg [7:0] dataMem_5_2__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_3__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_3__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_3__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_3__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_3__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_3__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_3__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_3__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_3__T_64_addr_pipe_0;
  reg  dataMem_5_3__T_167_en_pipe_0;
  reg [7:0] dataMem_5_3__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_4__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_4__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_4__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_4__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_4__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_4__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_4__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_4__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_4__T_64_addr_pipe_0;
  reg  dataMem_5_4__T_167_en_pipe_0;
  reg [7:0] dataMem_5_4__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_5__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_5__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_5__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_5__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_5__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_5__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_5__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_5__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_5__T_64_addr_pipe_0;
  reg  dataMem_5_5__T_167_en_pipe_0;
  reg [7:0] dataMem_5_5__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_6__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_6__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_6__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_6__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_6__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_6__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_6__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_6__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_6__T_64_addr_pipe_0;
  reg  dataMem_5_6__T_167_en_pipe_0;
  reg [7:0] dataMem_5_6__T_167_addr_pipe_0;
  reg [7:0] dataMem_5_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_7__T_64_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_7__T_64_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_7__T_167_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_7__T_167_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_7__T_376_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_5_7__T_376_addr; // @[AXICache.scala 721:45]
  wire  dataMem_5_7__T_376_mask; // @[AXICache.scala 721:45]
  wire  dataMem_5_7__T_376_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_5_7__T_64_addr_pipe_0;
  reg  dataMem_5_7__T_167_en_pipe_0;
  reg [7:0] dataMem_5_7__T_167_addr_pipe_0;
  reg [7:0] dataMem_6_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_0__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_0__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_0__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_0__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_0__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_0__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_0__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_0__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_0__T_74_addr_pipe_0;
  reg  dataMem_6_0__T_178_en_pipe_0;
  reg [7:0] dataMem_6_0__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_1__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_1__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_1__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_1__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_1__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_1__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_1__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_1__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_1__T_74_addr_pipe_0;
  reg  dataMem_6_1__T_178_en_pipe_0;
  reg [7:0] dataMem_6_1__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_2__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_2__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_2__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_2__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_2__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_2__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_2__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_2__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_2__T_74_addr_pipe_0;
  reg  dataMem_6_2__T_178_en_pipe_0;
  reg [7:0] dataMem_6_2__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_3__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_3__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_3__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_3__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_3__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_3__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_3__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_3__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_3__T_74_addr_pipe_0;
  reg  dataMem_6_3__T_178_en_pipe_0;
  reg [7:0] dataMem_6_3__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_4__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_4__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_4__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_4__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_4__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_4__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_4__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_4__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_4__T_74_addr_pipe_0;
  reg  dataMem_6_4__T_178_en_pipe_0;
  reg [7:0] dataMem_6_4__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_5__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_5__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_5__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_5__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_5__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_5__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_5__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_5__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_5__T_74_addr_pipe_0;
  reg  dataMem_6_5__T_178_en_pipe_0;
  reg [7:0] dataMem_6_5__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_6__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_6__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_6__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_6__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_6__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_6__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_6__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_6__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_6__T_74_addr_pipe_0;
  reg  dataMem_6_6__T_178_en_pipe_0;
  reg [7:0] dataMem_6_6__T_178_addr_pipe_0;
  reg [7:0] dataMem_6_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_7__T_74_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_7__T_74_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_7__T_178_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_7__T_178_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_7__T_395_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_6_7__T_395_addr; // @[AXICache.scala 721:45]
  wire  dataMem_6_7__T_395_mask; // @[AXICache.scala 721:45]
  wire  dataMem_6_7__T_395_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_6_7__T_74_addr_pipe_0;
  reg  dataMem_6_7__T_178_en_pipe_0;
  reg [7:0] dataMem_6_7__T_178_addr_pipe_0;
  reg [7:0] dataMem_7_0 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_0__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_0__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_0__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_0__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_0__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_0__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_0__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_0__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_0__T_84_addr_pipe_0;
  reg  dataMem_7_0__T_189_en_pipe_0;
  reg [7:0] dataMem_7_0__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_1 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_1__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_1__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_1__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_1__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_1__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_1__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_1__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_1__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_1__T_84_addr_pipe_0;
  reg  dataMem_7_1__T_189_en_pipe_0;
  reg [7:0] dataMem_7_1__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_2 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_2__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_2__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_2__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_2__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_2__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_2__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_2__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_2__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_2__T_84_addr_pipe_0;
  reg  dataMem_7_2__T_189_en_pipe_0;
  reg [7:0] dataMem_7_2__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_3 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_3__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_3__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_3__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_3__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_3__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_3__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_3__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_3__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_3__T_84_addr_pipe_0;
  reg  dataMem_7_3__T_189_en_pipe_0;
  reg [7:0] dataMem_7_3__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_4 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_4__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_4__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_4__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_4__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_4__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_4__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_4__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_4__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_4__T_84_addr_pipe_0;
  reg  dataMem_7_4__T_189_en_pipe_0;
  reg [7:0] dataMem_7_4__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_5 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_5__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_5__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_5__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_5__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_5__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_5__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_5__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_5__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_5__T_84_addr_pipe_0;
  reg  dataMem_7_5__T_189_en_pipe_0;
  reg [7:0] dataMem_7_5__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_6 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_6__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_6__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_6__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_6__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_6__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_6__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_6__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_6__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_6__T_84_addr_pipe_0;
  reg  dataMem_7_6__T_189_en_pipe_0;
  reg [7:0] dataMem_7_6__T_189_addr_pipe_0;
  reg [7:0] dataMem_7_7 [0:255]; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_7__T_84_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_7__T_84_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_7__T_189_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_7__T_189_addr; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_7__T_414_data; // @[AXICache.scala 721:45]
  wire [7:0] dataMem_7_7__T_414_addr; // @[AXICache.scala 721:45]
  wire  dataMem_7_7__T_414_mask; // @[AXICache.scala 721:45]
  wire  dataMem_7_7__T_414_en; // @[AXICache.scala 721:45]
  reg [7:0] dataMem_7_7__T_84_addr_pipe_0;
  reg  dataMem_7_7__T_189_en_pipe_0;
  reg [7:0] dataMem_7_7__T_189_addr_pipe_0;
  reg [2:0] state; // @[AXICache.scala 711:22]
  reg [2:0] flush_state; // @[AXICache.scala 714:28]
  reg  flush_mode; // @[AXICache.scala 715:27]
  reg [255:0] v; // @[AXICache.scala 718:18]
  reg [255:0] d; // @[AXICache.scala 719:18]
  reg [63:0] addr_reg; // @[AXICache.scala 723:21]
  reg [7:0] cpu_tag_reg; // @[AXICache.scala 724:24]
  reg [63:0] cpu_data; // @[AXICache.scala 726:21]
  reg [7:0] cpu_mask; // @[AXICache.scala 727:21]
  wire  _T = io_mem_rd_data_ready & io_mem_rd_data_valid; // @[Decoupled.scala 40:37]
  reg [2:0] read_count; // @[Counter.scala 29:33]
  wire  _T_1 = read_count == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_3 = read_count + 3'h1; // @[Counter.scala 39:22]
  wire  read_wrap_out = _T & _T_1; // @[Counter.scala 67:17]
  wire  _T_4 = io_mem_wr_data_ready & io_mem_wr_data_valid; // @[Decoupled.scala 40:37]
  reg [2:0] write_count; // @[Counter.scala 29:33]
  wire  _T_5 = write_count == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_7 = write_count + 3'h1; // @[Counter.scala 39:22]
  wire  write_wrap_out = _T_4 & _T_5; // @[Counter.scala 67:17]
  wire  _T_8 = flush_state == 3'h1; // @[AXICache.scala 734:51]
  reg [7:0] set_count; // @[Counter.scala 29:33]
  wire  _T_9 = set_count == 8'hff; // @[Counter.scala 38:24]
  wire [7:0] _T_11 = set_count + 8'h1; // @[Counter.scala 39:22]
  wire  set_wrap = _T_8 & _T_9; // @[Counter.scala 67:17]
  wire [7:0] _T_13 = set_count - 8'h1; // @[AXICache.scala 735:62]
  wire [63:0] _T_21 = {dataMem_0_7__T_14_data,dataMem_0_6__T_14_data,dataMem_0_5__T_14_data,dataMem_0_4__T_14_data,dataMem_0_3__T_14_data,dataMem_0_2__T_14_data,dataMem_0_1__T_14_data,dataMem_0_0__T_14_data}; // @[AXICache.scala 735:69]
  wire [63:0] _T_41 = {dataMem_2_7__T_34_data,dataMem_2_6__T_34_data,dataMem_2_5__T_34_data,dataMem_2_4__T_34_data,dataMem_2_3__T_34_data,dataMem_2_2__T_34_data,dataMem_2_1__T_34_data,dataMem_2_0__T_34_data}; // @[AXICache.scala 735:69]
  wire [63:0] _T_61 = {dataMem_4_7__T_54_data,dataMem_4_6__T_54_data,dataMem_4_5__T_54_data,dataMem_4_4__T_54_data,dataMem_4_3__T_54_data,dataMem_4_2__T_54_data,dataMem_4_1__T_54_data,dataMem_4_0__T_54_data}; // @[AXICache.scala 735:69]
  wire [63:0] _T_81 = {dataMem_6_7__T_74_data,dataMem_6_6__T_74_data,dataMem_6_5__T_74_data,dataMem_6_4__T_74_data,dataMem_6_3__T_74_data,dataMem_6_2__T_74_data,dataMem_6_1__T_74_data,dataMem_6_0__T_74_data}; // @[AXICache.scala 735:69]
  wire [127:0] _T_92 = {dataMem_1_7__T_24_data,dataMem_1_6__T_24_data,dataMem_1_5__T_24_data,dataMem_1_4__T_24_data,dataMem_1_3__T_24_data,dataMem_1_2__T_24_data,dataMem_1_1__T_24_data,dataMem_1_0__T_24_data,_T_21}; // @[Cat.scala 29:58]
  wire [255:0] _T_94 = {dataMem_3_7__T_44_data,dataMem_3_6__T_44_data,dataMem_3_5__T_44_data,dataMem_3_4__T_44_data,dataMem_3_3__T_44_data,dataMem_3_2__T_44_data,dataMem_3_1__T_44_data,dataMem_3_0__T_44_data,_T_41,_T_92}; // @[Cat.scala 29:58]
  wire [127:0] _T_95 = {dataMem_5_7__T_64_data,dataMem_5_6__T_64_data,dataMem_5_5__T_64_data,dataMem_5_4__T_64_data,dataMem_5_3__T_64_data,dataMem_5_2__T_64_data,dataMem_5_1__T_64_data,dataMem_5_0__T_64_data,_T_61}; // @[Cat.scala 29:58]
  wire [255:0] _T_97 = {dataMem_7_7__T_84_data,dataMem_7_6__T_84_data,dataMem_7_5__T_84_data,dataMem_7_4__T_84_data,dataMem_7_3__T_84_data,dataMem_7_2__T_84_data,dataMem_7_1__T_84_data,dataMem_7_0__T_84_data,_T_81,_T_95}; // @[Cat.scala 29:58]
  wire [511:0] dirty_cache_block = {_T_97,_T_94}; // @[Cat.scala 29:58]
  reg [49:0] block_rmeta_tag; // @[AXICache.scala 736:24]
  wire  is_idle = state == 3'h0; // @[AXICache.scala 740:23]
  wire  is_read = state == 3'h1; // @[AXICache.scala 741:23]
  wire  is_write = state == 3'h2; // @[AXICache.scala 742:24]
  wire  _T_98 = state == 3'h6; // @[AXICache.scala 743:24]
  wire  is_alloc = _T_98 & read_wrap_out; // @[AXICache.scala 743:37]
  reg  is_alloc_reg; // @[AXICache.scala 744:29]
  wire [7:0] idx_reg = addr_reg[13:6]; // @[AXICache.scala 754:25]
  wire [255:0] _T_211 = v >> idx_reg; // @[AXICache.scala 763:11]
  wire [49:0] tag_reg = addr_reg[63:14]; // @[AXICache.scala 753:25]
  wire  _T_213 = metaMem_tag_rmeta_data == tag_reg; // @[AXICache.scala 763:34]
  wire  hit = _T_211[0] & _T_213; // @[AXICache.scala 763:21]
  wire  _T_99 = hit | is_alloc_reg; // @[AXICache.scala 747:30]
  wire  _T_100 = is_write & _T_99; // @[AXICache.scala 747:22]
  wire  wen = _T_100 | is_alloc; // @[AXICache.scala 747:64]
  wire  _T_103 = ~wen; // @[AXICache.scala 748:13]
  wire  _T_104 = is_idle | is_read; // @[AXICache.scala 748:30]
  wire  _T_105 = _T_103 & _T_104; // @[AXICache.scala 748:18]
  reg  ren_reg; // @[AXICache.scala 749:24]
  wire [2:0] off_reg = addr_reg[5:3]; // @[AXICache.scala 755:25]
  wire [63:0] _T_119 = {dataMem_0_7__T_112_data,dataMem_0_6__T_112_data,dataMem_0_5__T_112_data,dataMem_0_4__T_112_data,dataMem_0_3__T_112_data,dataMem_0_2__T_112_data,dataMem_0_1__T_112_data,dataMem_0_0__T_112_data}; // @[AXICache.scala 758:50]
  wire [63:0] _T_141 = {dataMem_2_7__T_134_data,dataMem_2_6__T_134_data,dataMem_2_5__T_134_data,dataMem_2_4__T_134_data,dataMem_2_3__T_134_data,dataMem_2_2__T_134_data,dataMem_2_1__T_134_data,dataMem_2_0__T_134_data}; // @[AXICache.scala 758:50]
  wire [63:0] _T_163 = {dataMem_4_7__T_156_data,dataMem_4_6__T_156_data,dataMem_4_5__T_156_data,dataMem_4_4__T_156_data,dataMem_4_3__T_156_data,dataMem_4_2__T_156_data,dataMem_4_1__T_156_data,dataMem_4_0__T_156_data}; // @[AXICache.scala 758:50]
  wire [63:0] _T_185 = {dataMem_6_7__T_178_data,dataMem_6_6__T_178_data,dataMem_6_5__T_178_data,dataMem_6_4__T_178_data,dataMem_6_3__T_178_data,dataMem_6_2__T_178_data,dataMem_6_1__T_178_data,dataMem_6_0__T_178_data}; // @[AXICache.scala 758:50]
  wire [127:0] _T_197 = {dataMem_1_7__T_123_data,dataMem_1_6__T_123_data,dataMem_1_5__T_123_data,dataMem_1_4__T_123_data,dataMem_1_3__T_123_data,dataMem_1_2__T_123_data,dataMem_1_1__T_123_data,dataMem_1_0__T_123_data,_T_119}; // @[Cat.scala 29:58]
  wire [255:0] _T_199 = {dataMem_3_7__T_145_data,dataMem_3_6__T_145_data,dataMem_3_5__T_145_data,dataMem_3_4__T_145_data,dataMem_3_3__T_145_data,dataMem_3_2__T_145_data,dataMem_3_1__T_145_data,dataMem_3_0__T_145_data,_T_141,_T_197}; // @[Cat.scala 29:58]
  wire [127:0] _T_200 = {dataMem_5_7__T_167_data,dataMem_5_6__T_167_data,dataMem_5_5__T_167_data,dataMem_5_4__T_167_data,dataMem_5_3__T_167_data,dataMem_5_2__T_167_data,dataMem_5_1__T_167_data,dataMem_5_0__T_167_data,_T_163}; // @[Cat.scala 29:58]
  wire [255:0] _T_202 = {dataMem_7_7__T_189_data,dataMem_7_6__T_189_data,dataMem_7_5__T_189_data,dataMem_7_4__T_189_data,dataMem_7_3__T_189_data,dataMem_7_2__T_189_data,dataMem_7_1__T_189_data,dataMem_7_0__T_189_data,_T_185,_T_200}; // @[Cat.scala 29:58]
  wire [511:0] rdata = {_T_202,_T_199}; // @[Cat.scala 29:58]
  reg [511:0] rdata_buf; // @[Reg.scala 15:16]
  wire [511:0] _GEN_18 = ren_reg ? rdata : rdata_buf; // @[Reg.scala 16:19]
  reg [63:0] refill_buf_0; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_1; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_2; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_3; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_4; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_5; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_6; // @[AXICache.scala 760:23]
  reg [63:0] refill_buf_7; // @[AXICache.scala 760:23]
  wire [511:0] _T_209 = {refill_buf_7,refill_buf_6,refill_buf_5,refill_buf_4,refill_buf_3,refill_buf_2,refill_buf_1,refill_buf_0}; // @[AXICache.scala 761:43]
  wire [511:0] read = is_alloc_reg ? _T_209 : _GEN_18; // @[AXICache.scala 761:17]
  wire  _T_216 = is_read & hit; // @[AXICache.scala 765:58]
  wire  _T_217 = is_idle | _T_216; // @[AXICache.scala 765:31]
  wire [63:0] _GEN_20 = 3'h1 == off_reg ? read[127:64] : read[63:0]; // @[AXICache.scala 768:25]
  wire [63:0] _GEN_21 = 3'h2 == off_reg ? read[191:128] : _GEN_20; // @[AXICache.scala 768:25]
  wire [63:0] _GEN_22 = 3'h3 == off_reg ? read[255:192] : _GEN_21; // @[AXICache.scala 768:25]
  wire [63:0] _GEN_23 = 3'h4 == off_reg ? read[319:256] : _GEN_22; // @[AXICache.scala 768:25]
  wire [63:0] _GEN_24 = 3'h5 == off_reg ? read[383:320] : _GEN_23; // @[AXICache.scala 768:25]
  wire [63:0] _GEN_25 = 3'h6 == off_reg ? read[447:384] : _GEN_24; // @[AXICache.scala 768:25]
  wire  _T_229 = |cpu_mask; // @[AXICache.scala 769:79]
  wire  _T_230 = ~_T_229; // @[AXICache.scala 769:69]
  wire  _T_231 = is_alloc_reg & _T_230; // @[AXICache.scala 769:66]
  wire  _T_233 = io_cpu_req_ready & io_cpu_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_234 = ~is_alloc; // @[AXICache.scala 788:19]
  wire [5:0] _T_235 = {off_reg,3'h0}; // @[Cat.scala 29:58]
  wire [70:0] _GEN_407 = {{63'd0}, cpu_mask}; // @[AXICache.scala 788:40]
  wire [70:0] _T_236 = _GEN_407 << _T_235; // @[AXICache.scala 788:40]
  wire [71:0] _T_237 = {1'b0,$signed(_T_236)}; // @[AXICache.scala 788:91]
  wire [71:0] wmask = _T_234 ? $signed(_T_237) : $signed(-72'sh1); // @[AXICache.scala 788:18]
  wire [511:0] _T_241 = {cpu_data,cpu_data,cpu_data,cpu_data,cpu_data,cpu_data,cpu_data,cpu_data}; // @[Cat.scala 29:58]
  wire [511:0] _T_248 = {io_mem_rd_data_bits,refill_buf_6,refill_buf_5,refill_buf_4,refill_buf_3,refill_buf_2,refill_buf_1,refill_buf_0}; // @[Cat.scala 29:58]
  wire [511:0] wdata = _T_234 ? _T_241 : _T_248; // @[AXICache.scala 789:18]
  wire [255:0] _T_249 = 256'h1 << idx_reg; // @[AXICache.scala 793:18]
  wire [255:0] _T_250 = v | _T_249; // @[AXICache.scala 793:18]
  wire [255:0] _T_257 = d | _T_249; // @[AXICache.scala 794:18]
  wire [255:0] _T_258 = ~d; // @[AXICache.scala 794:18]
  wire [255:0] _T_259 = _T_258 | _T_249; // @[AXICache.scala 794:18]
  wire [255:0] _T_260 = ~_T_259; // @[AXICache.scala 794:18]
  wire [57:0] _T_415 = {tag_reg,idx_reg}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_408 = {_T_415, 6'h0}; // @[AXICache.scala 812:52]
  wire [64:0] _T_416 = {{1'd0}, _GEN_408}; // @[AXICache.scala 812:52]
  wire [255:0] _T_419 = v >> set_count; // @[AXICache.scala 823:25]
  wire [255:0] _T_421 = d >> set_count; // @[AXICache.scala 823:41]
  wire  is_block_dirty = _T_419[0] & _T_421[0]; // @[AXICache.scala 823:37]
  wire [57:0] _T_425 = {block_rmeta_tag,_T_13}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_409 = {_T_425, 6'h0}; // @[AXICache.scala 824:58]
  wire [64:0] block_addr = {{1'd0}, _GEN_409}; // @[AXICache.scala 824:58]
  wire [57:0] _T_432 = {metaMem_tag_rmeta_data,idx_reg}; // @[Cat.scala 29:58]
  wire [63:0] _GEN_410 = {_T_432, 6'h0}; // @[AXICache.scala 835:82]
  wire [64:0] _T_433 = {{1'd0}, _GEN_410}; // @[AXICache.scala 835:82]
  wire [64:0] _T_434 = flush_mode ? block_addr : _T_433; // @[AXICache.scala 835:33]
  wire [63:0] _GEN_324 = 3'h1 == write_count ? dirty_cache_block[127:64] : dirty_cache_block[63:0]; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_325 = 3'h2 == write_count ? dirty_cache_block[191:128] : _GEN_324; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_326 = 3'h3 == write_count ? dirty_cache_block[255:192] : _GEN_325; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_327 = 3'h4 == write_count ? dirty_cache_block[319:256] : _GEN_326; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_328 = 3'h5 == write_count ? dirty_cache_block[383:320] : _GEN_327; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_329 = 3'h6 == write_count ? dirty_cache_block[447:384] : _GEN_328; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_330 = 3'h7 == write_count ? dirty_cache_block[511:448] : _GEN_329; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_332 = 3'h1 == write_count ? read[127:64] : read[63:0]; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_333 = 3'h2 == write_count ? read[191:128] : _GEN_332; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_334 = 3'h3 == write_count ? read[255:192] : _GEN_333; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_335 = 3'h4 == write_count ? read[319:256] : _GEN_334; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_336 = 3'h5 == write_count ? read[383:320] : _GEN_335; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_337 = 3'h6 == write_count ? read[447:384] : _GEN_336; // @[AXICache.scala 840:29]
  wire [63:0] _GEN_338 = 3'h7 == write_count ? read[511:448] : _GEN_337; // @[AXICache.scala 840:29]
  wire [255:0] _T_456 = d >> idx_reg; // @[AXICache.scala 853:33]
  wire  is_dirty = _T_211[0] & _T_456[0]; // @[AXICache.scala 853:29]
  wire  _T_458 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_459 = |io_cpu_req_bits_mask; // @[AXICache.scala 857:43]
  wire  _T_461 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_464 = ~is_dirty; // @[AXICache.scala 869:32]
  wire  _T_465 = io_mem_wr_cmd_ready & io_mem_wr_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _T_466 = io_mem_rd_cmd_ready & io_mem_rd_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_344 = hit ? 1'h0 : is_dirty; // @[AXICache.scala 861:17]
  wire  _GEN_345 = hit ? 1'h0 : _T_464; // @[AXICache.scala 861:17]
  wire  _T_467 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_349 = _T_99 ? 1'h0 : is_dirty; // @[AXICache.scala 878:49]
  wire  _GEN_350 = _T_99 ? 1'h0 : _T_464; // @[AXICache.scala 878:49]
  wire  _T_473 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_474 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_475 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_477 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire  _GEN_359 = _T_474 ? 1'h0 : _T_475; // @[Conditional.scala 39:67]
  wire  _GEN_362 = _T_473 ? 1'h0 : _GEN_359; // @[Conditional.scala 39:67]
  wire  _GEN_364 = _T_467 & _GEN_349; // @[Conditional.scala 39:67]
  wire  _GEN_365 = _T_467 ? _GEN_350 : _GEN_362; // @[Conditional.scala 39:67]
  wire  _GEN_366 = _T_467 ? 1'h0 : _T_473; // @[Conditional.scala 39:67]
  wire  _GEN_368 = _T_461 ? _GEN_344 : _GEN_364; // @[Conditional.scala 39:67]
  wire  _GEN_369 = _T_461 ? _GEN_345 : _GEN_365; // @[Conditional.scala 39:67]
  wire  _GEN_370 = _T_461 ? 1'h0 : _GEN_366; // @[Conditional.scala 39:67]
  wire  _GEN_372 = _T_458 ? 1'h0 : _GEN_368; // @[Conditional.scala 40:58]
  wire  _GEN_373 = _T_458 ? 1'h0 : _GEN_369; // @[Conditional.scala 40:58]
  wire  _GEN_374 = _T_458 ? 1'h0 : _GEN_370; // @[Conditional.scala 40:58]
  wire  _T_480 = 3'h0 == flush_state; // @[Conditional.scala 37:30]
  wire  _GEN_376 = io_cpu_flush | flush_mode; // @[AXICache.scala 917:26]
  wire  _T_481 = 3'h1 == flush_state; // @[Conditional.scala 37:30]
  wire  _T_482 = 3'h2 == flush_state; // @[Conditional.scala 37:30]
  wire  _T_483 = 3'h3 == flush_state; // @[Conditional.scala 37:30]
  wire  _T_485 = 3'h4 == flush_state; // @[Conditional.scala 37:30]
  wire  _T_486 = 3'h5 == flush_state; // @[Conditional.scala 37:30]
  wire  _GEN_385 = _T_485 | _GEN_374; // @[Conditional.scala 39:67]
  wire  _GEN_387 = _T_483 | _GEN_372; // @[Conditional.scala 39:67]
  wire  _GEN_388 = _T_483 ? 1'h0 : _GEN_373; // @[Conditional.scala 39:67]
  wire  _GEN_390 = _T_483 ? _GEN_374 : _GEN_385; // @[Conditional.scala 39:67]
  wire  _GEN_392 = _T_482 ? _GEN_372 : _GEN_387; // @[Conditional.scala 39:67]
  wire  _GEN_393 = _T_482 ? _GEN_373 : _GEN_388; // @[Conditional.scala 39:67]
  wire  _GEN_394 = _T_482 ? _GEN_374 : _GEN_390; // @[Conditional.scala 39:67]
  wire  _GEN_395 = _T_481 & set_wrap; // @[Conditional.scala 39:67]
  wire  _GEN_398 = _T_481 ? _GEN_372 : _GEN_392; // @[Conditional.scala 39:67]
  wire  _GEN_399 = _T_481 ? _GEN_373 : _GEN_393; // @[Conditional.scala 39:67]
  wire  _GEN_400 = _T_481 ? _GEN_374 : _GEN_394; // @[Conditional.scala 39:67]
  assign metaMem_tag_rmeta_addr = metaMem_tag_rmeta_addr_pipe_0;
  assign metaMem_tag_rmeta_data = metaMem_tag[metaMem_tag_rmeta_addr]; // @[AXICache.scala 720:28]
  assign metaMem_tag__T_431_addr = metaMem_tag__T_431_addr_pipe_0;
  assign metaMem_tag__T_431_data = metaMem_tag[metaMem_tag__T_431_addr]; // @[AXICache.scala 720:28]
  assign metaMem_tag__T_262_data = addr_reg[63:14];
  assign metaMem_tag__T_262_addr = addr_reg[13:6];
  assign metaMem_tag__T_262_mask = 1'h1;
  assign metaMem_tag__T_262_en = wen & is_alloc;
  assign dataMem_0_0__T_14_addr = dataMem_0_0__T_14_addr_pipe_0;
  assign dataMem_0_0__T_14_data = dataMem_0_0[dataMem_0_0__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_0__T_112_addr = dataMem_0_0__T_112_addr_pipe_0;
  assign dataMem_0_0__T_112_data = dataMem_0_0[dataMem_0_0__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_0__T_281_data = wdata[7:0];
  assign dataMem_0_0__T_281_addr = addr_reg[13:6];
  assign dataMem_0_0__T_281_mask = wmask[0];
  assign dataMem_0_0__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_1__T_14_addr = dataMem_0_1__T_14_addr_pipe_0;
  assign dataMem_0_1__T_14_data = dataMem_0_1[dataMem_0_1__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_1__T_112_addr = dataMem_0_1__T_112_addr_pipe_0;
  assign dataMem_0_1__T_112_data = dataMem_0_1[dataMem_0_1__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_1__T_281_data = wdata[15:8];
  assign dataMem_0_1__T_281_addr = addr_reg[13:6];
  assign dataMem_0_1__T_281_mask = wmask[1];
  assign dataMem_0_1__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_2__T_14_addr = dataMem_0_2__T_14_addr_pipe_0;
  assign dataMem_0_2__T_14_data = dataMem_0_2[dataMem_0_2__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_2__T_112_addr = dataMem_0_2__T_112_addr_pipe_0;
  assign dataMem_0_2__T_112_data = dataMem_0_2[dataMem_0_2__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_2__T_281_data = wdata[23:16];
  assign dataMem_0_2__T_281_addr = addr_reg[13:6];
  assign dataMem_0_2__T_281_mask = wmask[2];
  assign dataMem_0_2__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_3__T_14_addr = dataMem_0_3__T_14_addr_pipe_0;
  assign dataMem_0_3__T_14_data = dataMem_0_3[dataMem_0_3__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_3__T_112_addr = dataMem_0_3__T_112_addr_pipe_0;
  assign dataMem_0_3__T_112_data = dataMem_0_3[dataMem_0_3__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_3__T_281_data = wdata[31:24];
  assign dataMem_0_3__T_281_addr = addr_reg[13:6];
  assign dataMem_0_3__T_281_mask = wmask[3];
  assign dataMem_0_3__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_4__T_14_addr = dataMem_0_4__T_14_addr_pipe_0;
  assign dataMem_0_4__T_14_data = dataMem_0_4[dataMem_0_4__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_4__T_112_addr = dataMem_0_4__T_112_addr_pipe_0;
  assign dataMem_0_4__T_112_data = dataMem_0_4[dataMem_0_4__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_4__T_281_data = wdata[39:32];
  assign dataMem_0_4__T_281_addr = addr_reg[13:6];
  assign dataMem_0_4__T_281_mask = wmask[4];
  assign dataMem_0_4__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_5__T_14_addr = dataMem_0_5__T_14_addr_pipe_0;
  assign dataMem_0_5__T_14_data = dataMem_0_5[dataMem_0_5__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_5__T_112_addr = dataMem_0_5__T_112_addr_pipe_0;
  assign dataMem_0_5__T_112_data = dataMem_0_5[dataMem_0_5__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_5__T_281_data = wdata[47:40];
  assign dataMem_0_5__T_281_addr = addr_reg[13:6];
  assign dataMem_0_5__T_281_mask = wmask[5];
  assign dataMem_0_5__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_6__T_14_addr = dataMem_0_6__T_14_addr_pipe_0;
  assign dataMem_0_6__T_14_data = dataMem_0_6[dataMem_0_6__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_6__T_112_addr = dataMem_0_6__T_112_addr_pipe_0;
  assign dataMem_0_6__T_112_data = dataMem_0_6[dataMem_0_6__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_6__T_281_data = wdata[55:48];
  assign dataMem_0_6__T_281_addr = addr_reg[13:6];
  assign dataMem_0_6__T_281_mask = wmask[6];
  assign dataMem_0_6__T_281_en = _T_100 | is_alloc;
  assign dataMem_0_7__T_14_addr = dataMem_0_7__T_14_addr_pipe_0;
  assign dataMem_0_7__T_14_data = dataMem_0_7[dataMem_0_7__T_14_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_7__T_112_addr = dataMem_0_7__T_112_addr_pipe_0;
  assign dataMem_0_7__T_112_data = dataMem_0_7[dataMem_0_7__T_112_addr]; // @[AXICache.scala 721:45]
  assign dataMem_0_7__T_281_data = wdata[63:56];
  assign dataMem_0_7__T_281_addr = addr_reg[13:6];
  assign dataMem_0_7__T_281_mask = wmask[7];
  assign dataMem_0_7__T_281_en = _T_100 | is_alloc;
  assign dataMem_1_0__T_24_addr = dataMem_1_0__T_24_addr_pipe_0;
  assign dataMem_1_0__T_24_data = dataMem_1_0[dataMem_1_0__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_0__T_123_addr = dataMem_1_0__T_123_addr_pipe_0;
  assign dataMem_1_0__T_123_data = dataMem_1_0[dataMem_1_0__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_0__T_300_data = wdata[71:64];
  assign dataMem_1_0__T_300_addr = addr_reg[13:6];
  assign dataMem_1_0__T_300_mask = wmask[8];
  assign dataMem_1_0__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_1__T_24_addr = dataMem_1_1__T_24_addr_pipe_0;
  assign dataMem_1_1__T_24_data = dataMem_1_1[dataMem_1_1__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_1__T_123_addr = dataMem_1_1__T_123_addr_pipe_0;
  assign dataMem_1_1__T_123_data = dataMem_1_1[dataMem_1_1__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_1__T_300_data = wdata[79:72];
  assign dataMem_1_1__T_300_addr = addr_reg[13:6];
  assign dataMem_1_1__T_300_mask = wmask[9];
  assign dataMem_1_1__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_2__T_24_addr = dataMem_1_2__T_24_addr_pipe_0;
  assign dataMem_1_2__T_24_data = dataMem_1_2[dataMem_1_2__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_2__T_123_addr = dataMem_1_2__T_123_addr_pipe_0;
  assign dataMem_1_2__T_123_data = dataMem_1_2[dataMem_1_2__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_2__T_300_data = wdata[87:80];
  assign dataMem_1_2__T_300_addr = addr_reg[13:6];
  assign dataMem_1_2__T_300_mask = wmask[10];
  assign dataMem_1_2__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_3__T_24_addr = dataMem_1_3__T_24_addr_pipe_0;
  assign dataMem_1_3__T_24_data = dataMem_1_3[dataMem_1_3__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_3__T_123_addr = dataMem_1_3__T_123_addr_pipe_0;
  assign dataMem_1_3__T_123_data = dataMem_1_3[dataMem_1_3__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_3__T_300_data = wdata[95:88];
  assign dataMem_1_3__T_300_addr = addr_reg[13:6];
  assign dataMem_1_3__T_300_mask = wmask[11];
  assign dataMem_1_3__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_4__T_24_addr = dataMem_1_4__T_24_addr_pipe_0;
  assign dataMem_1_4__T_24_data = dataMem_1_4[dataMem_1_4__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_4__T_123_addr = dataMem_1_4__T_123_addr_pipe_0;
  assign dataMem_1_4__T_123_data = dataMem_1_4[dataMem_1_4__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_4__T_300_data = wdata[103:96];
  assign dataMem_1_4__T_300_addr = addr_reg[13:6];
  assign dataMem_1_4__T_300_mask = wmask[12];
  assign dataMem_1_4__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_5__T_24_addr = dataMem_1_5__T_24_addr_pipe_0;
  assign dataMem_1_5__T_24_data = dataMem_1_5[dataMem_1_5__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_5__T_123_addr = dataMem_1_5__T_123_addr_pipe_0;
  assign dataMem_1_5__T_123_data = dataMem_1_5[dataMem_1_5__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_5__T_300_data = wdata[111:104];
  assign dataMem_1_5__T_300_addr = addr_reg[13:6];
  assign dataMem_1_5__T_300_mask = wmask[13];
  assign dataMem_1_5__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_6__T_24_addr = dataMem_1_6__T_24_addr_pipe_0;
  assign dataMem_1_6__T_24_data = dataMem_1_6[dataMem_1_6__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_6__T_123_addr = dataMem_1_6__T_123_addr_pipe_0;
  assign dataMem_1_6__T_123_data = dataMem_1_6[dataMem_1_6__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_6__T_300_data = wdata[119:112];
  assign dataMem_1_6__T_300_addr = addr_reg[13:6];
  assign dataMem_1_6__T_300_mask = wmask[14];
  assign dataMem_1_6__T_300_en = _T_100 | is_alloc;
  assign dataMem_1_7__T_24_addr = dataMem_1_7__T_24_addr_pipe_0;
  assign dataMem_1_7__T_24_data = dataMem_1_7[dataMem_1_7__T_24_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_7__T_123_addr = dataMem_1_7__T_123_addr_pipe_0;
  assign dataMem_1_7__T_123_data = dataMem_1_7[dataMem_1_7__T_123_addr]; // @[AXICache.scala 721:45]
  assign dataMem_1_7__T_300_data = wdata[127:120];
  assign dataMem_1_7__T_300_addr = addr_reg[13:6];
  assign dataMem_1_7__T_300_mask = wmask[15];
  assign dataMem_1_7__T_300_en = _T_100 | is_alloc;
  assign dataMem_2_0__T_34_addr = dataMem_2_0__T_34_addr_pipe_0;
  assign dataMem_2_0__T_34_data = dataMem_2_0[dataMem_2_0__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_0__T_134_addr = dataMem_2_0__T_134_addr_pipe_0;
  assign dataMem_2_0__T_134_data = dataMem_2_0[dataMem_2_0__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_0__T_319_data = wdata[135:128];
  assign dataMem_2_0__T_319_addr = addr_reg[13:6];
  assign dataMem_2_0__T_319_mask = wmask[16];
  assign dataMem_2_0__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_1__T_34_addr = dataMem_2_1__T_34_addr_pipe_0;
  assign dataMem_2_1__T_34_data = dataMem_2_1[dataMem_2_1__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_1__T_134_addr = dataMem_2_1__T_134_addr_pipe_0;
  assign dataMem_2_1__T_134_data = dataMem_2_1[dataMem_2_1__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_1__T_319_data = wdata[143:136];
  assign dataMem_2_1__T_319_addr = addr_reg[13:6];
  assign dataMem_2_1__T_319_mask = wmask[17];
  assign dataMem_2_1__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_2__T_34_addr = dataMem_2_2__T_34_addr_pipe_0;
  assign dataMem_2_2__T_34_data = dataMem_2_2[dataMem_2_2__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_2__T_134_addr = dataMem_2_2__T_134_addr_pipe_0;
  assign dataMem_2_2__T_134_data = dataMem_2_2[dataMem_2_2__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_2__T_319_data = wdata[151:144];
  assign dataMem_2_2__T_319_addr = addr_reg[13:6];
  assign dataMem_2_2__T_319_mask = wmask[18];
  assign dataMem_2_2__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_3__T_34_addr = dataMem_2_3__T_34_addr_pipe_0;
  assign dataMem_2_3__T_34_data = dataMem_2_3[dataMem_2_3__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_3__T_134_addr = dataMem_2_3__T_134_addr_pipe_0;
  assign dataMem_2_3__T_134_data = dataMem_2_3[dataMem_2_3__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_3__T_319_data = wdata[159:152];
  assign dataMem_2_3__T_319_addr = addr_reg[13:6];
  assign dataMem_2_3__T_319_mask = wmask[19];
  assign dataMem_2_3__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_4__T_34_addr = dataMem_2_4__T_34_addr_pipe_0;
  assign dataMem_2_4__T_34_data = dataMem_2_4[dataMem_2_4__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_4__T_134_addr = dataMem_2_4__T_134_addr_pipe_0;
  assign dataMem_2_4__T_134_data = dataMem_2_4[dataMem_2_4__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_4__T_319_data = wdata[167:160];
  assign dataMem_2_4__T_319_addr = addr_reg[13:6];
  assign dataMem_2_4__T_319_mask = wmask[20];
  assign dataMem_2_4__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_5__T_34_addr = dataMem_2_5__T_34_addr_pipe_0;
  assign dataMem_2_5__T_34_data = dataMem_2_5[dataMem_2_5__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_5__T_134_addr = dataMem_2_5__T_134_addr_pipe_0;
  assign dataMem_2_5__T_134_data = dataMem_2_5[dataMem_2_5__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_5__T_319_data = wdata[175:168];
  assign dataMem_2_5__T_319_addr = addr_reg[13:6];
  assign dataMem_2_5__T_319_mask = wmask[21];
  assign dataMem_2_5__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_6__T_34_addr = dataMem_2_6__T_34_addr_pipe_0;
  assign dataMem_2_6__T_34_data = dataMem_2_6[dataMem_2_6__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_6__T_134_addr = dataMem_2_6__T_134_addr_pipe_0;
  assign dataMem_2_6__T_134_data = dataMem_2_6[dataMem_2_6__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_6__T_319_data = wdata[183:176];
  assign dataMem_2_6__T_319_addr = addr_reg[13:6];
  assign dataMem_2_6__T_319_mask = wmask[22];
  assign dataMem_2_6__T_319_en = _T_100 | is_alloc;
  assign dataMem_2_7__T_34_addr = dataMem_2_7__T_34_addr_pipe_0;
  assign dataMem_2_7__T_34_data = dataMem_2_7[dataMem_2_7__T_34_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_7__T_134_addr = dataMem_2_7__T_134_addr_pipe_0;
  assign dataMem_2_7__T_134_data = dataMem_2_7[dataMem_2_7__T_134_addr]; // @[AXICache.scala 721:45]
  assign dataMem_2_7__T_319_data = wdata[191:184];
  assign dataMem_2_7__T_319_addr = addr_reg[13:6];
  assign dataMem_2_7__T_319_mask = wmask[23];
  assign dataMem_2_7__T_319_en = _T_100 | is_alloc;
  assign dataMem_3_0__T_44_addr = dataMem_3_0__T_44_addr_pipe_0;
  assign dataMem_3_0__T_44_data = dataMem_3_0[dataMem_3_0__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_0__T_145_addr = dataMem_3_0__T_145_addr_pipe_0;
  assign dataMem_3_0__T_145_data = dataMem_3_0[dataMem_3_0__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_0__T_338_data = wdata[199:192];
  assign dataMem_3_0__T_338_addr = addr_reg[13:6];
  assign dataMem_3_0__T_338_mask = wmask[24];
  assign dataMem_3_0__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_1__T_44_addr = dataMem_3_1__T_44_addr_pipe_0;
  assign dataMem_3_1__T_44_data = dataMem_3_1[dataMem_3_1__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_1__T_145_addr = dataMem_3_1__T_145_addr_pipe_0;
  assign dataMem_3_1__T_145_data = dataMem_3_1[dataMem_3_1__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_1__T_338_data = wdata[207:200];
  assign dataMem_3_1__T_338_addr = addr_reg[13:6];
  assign dataMem_3_1__T_338_mask = wmask[25];
  assign dataMem_3_1__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_2__T_44_addr = dataMem_3_2__T_44_addr_pipe_0;
  assign dataMem_3_2__T_44_data = dataMem_3_2[dataMem_3_2__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_2__T_145_addr = dataMem_3_2__T_145_addr_pipe_0;
  assign dataMem_3_2__T_145_data = dataMem_3_2[dataMem_3_2__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_2__T_338_data = wdata[215:208];
  assign dataMem_3_2__T_338_addr = addr_reg[13:6];
  assign dataMem_3_2__T_338_mask = wmask[26];
  assign dataMem_3_2__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_3__T_44_addr = dataMem_3_3__T_44_addr_pipe_0;
  assign dataMem_3_3__T_44_data = dataMem_3_3[dataMem_3_3__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_3__T_145_addr = dataMem_3_3__T_145_addr_pipe_0;
  assign dataMem_3_3__T_145_data = dataMem_3_3[dataMem_3_3__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_3__T_338_data = wdata[223:216];
  assign dataMem_3_3__T_338_addr = addr_reg[13:6];
  assign dataMem_3_3__T_338_mask = wmask[27];
  assign dataMem_3_3__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_4__T_44_addr = dataMem_3_4__T_44_addr_pipe_0;
  assign dataMem_3_4__T_44_data = dataMem_3_4[dataMem_3_4__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_4__T_145_addr = dataMem_3_4__T_145_addr_pipe_0;
  assign dataMem_3_4__T_145_data = dataMem_3_4[dataMem_3_4__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_4__T_338_data = wdata[231:224];
  assign dataMem_3_4__T_338_addr = addr_reg[13:6];
  assign dataMem_3_4__T_338_mask = wmask[28];
  assign dataMem_3_4__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_5__T_44_addr = dataMem_3_5__T_44_addr_pipe_0;
  assign dataMem_3_5__T_44_data = dataMem_3_5[dataMem_3_5__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_5__T_145_addr = dataMem_3_5__T_145_addr_pipe_0;
  assign dataMem_3_5__T_145_data = dataMem_3_5[dataMem_3_5__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_5__T_338_data = wdata[239:232];
  assign dataMem_3_5__T_338_addr = addr_reg[13:6];
  assign dataMem_3_5__T_338_mask = wmask[29];
  assign dataMem_3_5__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_6__T_44_addr = dataMem_3_6__T_44_addr_pipe_0;
  assign dataMem_3_6__T_44_data = dataMem_3_6[dataMem_3_6__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_6__T_145_addr = dataMem_3_6__T_145_addr_pipe_0;
  assign dataMem_3_6__T_145_data = dataMem_3_6[dataMem_3_6__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_6__T_338_data = wdata[247:240];
  assign dataMem_3_6__T_338_addr = addr_reg[13:6];
  assign dataMem_3_6__T_338_mask = wmask[30];
  assign dataMem_3_6__T_338_en = _T_100 | is_alloc;
  assign dataMem_3_7__T_44_addr = dataMem_3_7__T_44_addr_pipe_0;
  assign dataMem_3_7__T_44_data = dataMem_3_7[dataMem_3_7__T_44_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_7__T_145_addr = dataMem_3_7__T_145_addr_pipe_0;
  assign dataMem_3_7__T_145_data = dataMem_3_7[dataMem_3_7__T_145_addr]; // @[AXICache.scala 721:45]
  assign dataMem_3_7__T_338_data = wdata[255:248];
  assign dataMem_3_7__T_338_addr = addr_reg[13:6];
  assign dataMem_3_7__T_338_mask = wmask[31];
  assign dataMem_3_7__T_338_en = _T_100 | is_alloc;
  assign dataMem_4_0__T_54_addr = dataMem_4_0__T_54_addr_pipe_0;
  assign dataMem_4_0__T_54_data = dataMem_4_0[dataMem_4_0__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_0__T_156_addr = dataMem_4_0__T_156_addr_pipe_0;
  assign dataMem_4_0__T_156_data = dataMem_4_0[dataMem_4_0__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_0__T_357_data = wdata[263:256];
  assign dataMem_4_0__T_357_addr = addr_reg[13:6];
  assign dataMem_4_0__T_357_mask = wmask[32];
  assign dataMem_4_0__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_1__T_54_addr = dataMem_4_1__T_54_addr_pipe_0;
  assign dataMem_4_1__T_54_data = dataMem_4_1[dataMem_4_1__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_1__T_156_addr = dataMem_4_1__T_156_addr_pipe_0;
  assign dataMem_4_1__T_156_data = dataMem_4_1[dataMem_4_1__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_1__T_357_data = wdata[271:264];
  assign dataMem_4_1__T_357_addr = addr_reg[13:6];
  assign dataMem_4_1__T_357_mask = wmask[33];
  assign dataMem_4_1__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_2__T_54_addr = dataMem_4_2__T_54_addr_pipe_0;
  assign dataMem_4_2__T_54_data = dataMem_4_2[dataMem_4_2__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_2__T_156_addr = dataMem_4_2__T_156_addr_pipe_0;
  assign dataMem_4_2__T_156_data = dataMem_4_2[dataMem_4_2__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_2__T_357_data = wdata[279:272];
  assign dataMem_4_2__T_357_addr = addr_reg[13:6];
  assign dataMem_4_2__T_357_mask = wmask[34];
  assign dataMem_4_2__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_3__T_54_addr = dataMem_4_3__T_54_addr_pipe_0;
  assign dataMem_4_3__T_54_data = dataMem_4_3[dataMem_4_3__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_3__T_156_addr = dataMem_4_3__T_156_addr_pipe_0;
  assign dataMem_4_3__T_156_data = dataMem_4_3[dataMem_4_3__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_3__T_357_data = wdata[287:280];
  assign dataMem_4_3__T_357_addr = addr_reg[13:6];
  assign dataMem_4_3__T_357_mask = wmask[35];
  assign dataMem_4_3__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_4__T_54_addr = dataMem_4_4__T_54_addr_pipe_0;
  assign dataMem_4_4__T_54_data = dataMem_4_4[dataMem_4_4__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_4__T_156_addr = dataMem_4_4__T_156_addr_pipe_0;
  assign dataMem_4_4__T_156_data = dataMem_4_4[dataMem_4_4__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_4__T_357_data = wdata[295:288];
  assign dataMem_4_4__T_357_addr = addr_reg[13:6];
  assign dataMem_4_4__T_357_mask = wmask[36];
  assign dataMem_4_4__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_5__T_54_addr = dataMem_4_5__T_54_addr_pipe_0;
  assign dataMem_4_5__T_54_data = dataMem_4_5[dataMem_4_5__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_5__T_156_addr = dataMem_4_5__T_156_addr_pipe_0;
  assign dataMem_4_5__T_156_data = dataMem_4_5[dataMem_4_5__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_5__T_357_data = wdata[303:296];
  assign dataMem_4_5__T_357_addr = addr_reg[13:6];
  assign dataMem_4_5__T_357_mask = wmask[37];
  assign dataMem_4_5__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_6__T_54_addr = dataMem_4_6__T_54_addr_pipe_0;
  assign dataMem_4_6__T_54_data = dataMem_4_6[dataMem_4_6__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_6__T_156_addr = dataMem_4_6__T_156_addr_pipe_0;
  assign dataMem_4_6__T_156_data = dataMem_4_6[dataMem_4_6__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_6__T_357_data = wdata[311:304];
  assign dataMem_4_6__T_357_addr = addr_reg[13:6];
  assign dataMem_4_6__T_357_mask = wmask[38];
  assign dataMem_4_6__T_357_en = _T_100 | is_alloc;
  assign dataMem_4_7__T_54_addr = dataMem_4_7__T_54_addr_pipe_0;
  assign dataMem_4_7__T_54_data = dataMem_4_7[dataMem_4_7__T_54_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_7__T_156_addr = dataMem_4_7__T_156_addr_pipe_0;
  assign dataMem_4_7__T_156_data = dataMem_4_7[dataMem_4_7__T_156_addr]; // @[AXICache.scala 721:45]
  assign dataMem_4_7__T_357_data = wdata[319:312];
  assign dataMem_4_7__T_357_addr = addr_reg[13:6];
  assign dataMem_4_7__T_357_mask = wmask[39];
  assign dataMem_4_7__T_357_en = _T_100 | is_alloc;
  assign dataMem_5_0__T_64_addr = dataMem_5_0__T_64_addr_pipe_0;
  assign dataMem_5_0__T_64_data = dataMem_5_0[dataMem_5_0__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_0__T_167_addr = dataMem_5_0__T_167_addr_pipe_0;
  assign dataMem_5_0__T_167_data = dataMem_5_0[dataMem_5_0__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_0__T_376_data = wdata[327:320];
  assign dataMem_5_0__T_376_addr = addr_reg[13:6];
  assign dataMem_5_0__T_376_mask = wmask[40];
  assign dataMem_5_0__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_1__T_64_addr = dataMem_5_1__T_64_addr_pipe_0;
  assign dataMem_5_1__T_64_data = dataMem_5_1[dataMem_5_1__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_1__T_167_addr = dataMem_5_1__T_167_addr_pipe_0;
  assign dataMem_5_1__T_167_data = dataMem_5_1[dataMem_5_1__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_1__T_376_data = wdata[335:328];
  assign dataMem_5_1__T_376_addr = addr_reg[13:6];
  assign dataMem_5_1__T_376_mask = wmask[41];
  assign dataMem_5_1__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_2__T_64_addr = dataMem_5_2__T_64_addr_pipe_0;
  assign dataMem_5_2__T_64_data = dataMem_5_2[dataMem_5_2__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_2__T_167_addr = dataMem_5_2__T_167_addr_pipe_0;
  assign dataMem_5_2__T_167_data = dataMem_5_2[dataMem_5_2__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_2__T_376_data = wdata[343:336];
  assign dataMem_5_2__T_376_addr = addr_reg[13:6];
  assign dataMem_5_2__T_376_mask = wmask[42];
  assign dataMem_5_2__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_3__T_64_addr = dataMem_5_3__T_64_addr_pipe_0;
  assign dataMem_5_3__T_64_data = dataMem_5_3[dataMem_5_3__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_3__T_167_addr = dataMem_5_3__T_167_addr_pipe_0;
  assign dataMem_5_3__T_167_data = dataMem_5_3[dataMem_5_3__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_3__T_376_data = wdata[351:344];
  assign dataMem_5_3__T_376_addr = addr_reg[13:6];
  assign dataMem_5_3__T_376_mask = wmask[43];
  assign dataMem_5_3__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_4__T_64_addr = dataMem_5_4__T_64_addr_pipe_0;
  assign dataMem_5_4__T_64_data = dataMem_5_4[dataMem_5_4__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_4__T_167_addr = dataMem_5_4__T_167_addr_pipe_0;
  assign dataMem_5_4__T_167_data = dataMem_5_4[dataMem_5_4__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_4__T_376_data = wdata[359:352];
  assign dataMem_5_4__T_376_addr = addr_reg[13:6];
  assign dataMem_5_4__T_376_mask = wmask[44];
  assign dataMem_5_4__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_5__T_64_addr = dataMem_5_5__T_64_addr_pipe_0;
  assign dataMem_5_5__T_64_data = dataMem_5_5[dataMem_5_5__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_5__T_167_addr = dataMem_5_5__T_167_addr_pipe_0;
  assign dataMem_5_5__T_167_data = dataMem_5_5[dataMem_5_5__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_5__T_376_data = wdata[367:360];
  assign dataMem_5_5__T_376_addr = addr_reg[13:6];
  assign dataMem_5_5__T_376_mask = wmask[45];
  assign dataMem_5_5__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_6__T_64_addr = dataMem_5_6__T_64_addr_pipe_0;
  assign dataMem_5_6__T_64_data = dataMem_5_6[dataMem_5_6__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_6__T_167_addr = dataMem_5_6__T_167_addr_pipe_0;
  assign dataMem_5_6__T_167_data = dataMem_5_6[dataMem_5_6__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_6__T_376_data = wdata[375:368];
  assign dataMem_5_6__T_376_addr = addr_reg[13:6];
  assign dataMem_5_6__T_376_mask = wmask[46];
  assign dataMem_5_6__T_376_en = _T_100 | is_alloc;
  assign dataMem_5_7__T_64_addr = dataMem_5_7__T_64_addr_pipe_0;
  assign dataMem_5_7__T_64_data = dataMem_5_7[dataMem_5_7__T_64_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_7__T_167_addr = dataMem_5_7__T_167_addr_pipe_0;
  assign dataMem_5_7__T_167_data = dataMem_5_7[dataMem_5_7__T_167_addr]; // @[AXICache.scala 721:45]
  assign dataMem_5_7__T_376_data = wdata[383:376];
  assign dataMem_5_7__T_376_addr = addr_reg[13:6];
  assign dataMem_5_7__T_376_mask = wmask[47];
  assign dataMem_5_7__T_376_en = _T_100 | is_alloc;
  assign dataMem_6_0__T_74_addr = dataMem_6_0__T_74_addr_pipe_0;
  assign dataMem_6_0__T_74_data = dataMem_6_0[dataMem_6_0__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_0__T_178_addr = dataMem_6_0__T_178_addr_pipe_0;
  assign dataMem_6_0__T_178_data = dataMem_6_0[dataMem_6_0__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_0__T_395_data = wdata[391:384];
  assign dataMem_6_0__T_395_addr = addr_reg[13:6];
  assign dataMem_6_0__T_395_mask = wmask[48];
  assign dataMem_6_0__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_1__T_74_addr = dataMem_6_1__T_74_addr_pipe_0;
  assign dataMem_6_1__T_74_data = dataMem_6_1[dataMem_6_1__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_1__T_178_addr = dataMem_6_1__T_178_addr_pipe_0;
  assign dataMem_6_1__T_178_data = dataMem_6_1[dataMem_6_1__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_1__T_395_data = wdata[399:392];
  assign dataMem_6_1__T_395_addr = addr_reg[13:6];
  assign dataMem_6_1__T_395_mask = wmask[49];
  assign dataMem_6_1__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_2__T_74_addr = dataMem_6_2__T_74_addr_pipe_0;
  assign dataMem_6_2__T_74_data = dataMem_6_2[dataMem_6_2__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_2__T_178_addr = dataMem_6_2__T_178_addr_pipe_0;
  assign dataMem_6_2__T_178_data = dataMem_6_2[dataMem_6_2__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_2__T_395_data = wdata[407:400];
  assign dataMem_6_2__T_395_addr = addr_reg[13:6];
  assign dataMem_6_2__T_395_mask = wmask[50];
  assign dataMem_6_2__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_3__T_74_addr = dataMem_6_3__T_74_addr_pipe_0;
  assign dataMem_6_3__T_74_data = dataMem_6_3[dataMem_6_3__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_3__T_178_addr = dataMem_6_3__T_178_addr_pipe_0;
  assign dataMem_6_3__T_178_data = dataMem_6_3[dataMem_6_3__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_3__T_395_data = wdata[415:408];
  assign dataMem_6_3__T_395_addr = addr_reg[13:6];
  assign dataMem_6_3__T_395_mask = wmask[51];
  assign dataMem_6_3__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_4__T_74_addr = dataMem_6_4__T_74_addr_pipe_0;
  assign dataMem_6_4__T_74_data = dataMem_6_4[dataMem_6_4__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_4__T_178_addr = dataMem_6_4__T_178_addr_pipe_0;
  assign dataMem_6_4__T_178_data = dataMem_6_4[dataMem_6_4__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_4__T_395_data = wdata[423:416];
  assign dataMem_6_4__T_395_addr = addr_reg[13:6];
  assign dataMem_6_4__T_395_mask = wmask[52];
  assign dataMem_6_4__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_5__T_74_addr = dataMem_6_5__T_74_addr_pipe_0;
  assign dataMem_6_5__T_74_data = dataMem_6_5[dataMem_6_5__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_5__T_178_addr = dataMem_6_5__T_178_addr_pipe_0;
  assign dataMem_6_5__T_178_data = dataMem_6_5[dataMem_6_5__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_5__T_395_data = wdata[431:424];
  assign dataMem_6_5__T_395_addr = addr_reg[13:6];
  assign dataMem_6_5__T_395_mask = wmask[53];
  assign dataMem_6_5__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_6__T_74_addr = dataMem_6_6__T_74_addr_pipe_0;
  assign dataMem_6_6__T_74_data = dataMem_6_6[dataMem_6_6__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_6__T_178_addr = dataMem_6_6__T_178_addr_pipe_0;
  assign dataMem_6_6__T_178_data = dataMem_6_6[dataMem_6_6__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_6__T_395_data = wdata[439:432];
  assign dataMem_6_6__T_395_addr = addr_reg[13:6];
  assign dataMem_6_6__T_395_mask = wmask[54];
  assign dataMem_6_6__T_395_en = _T_100 | is_alloc;
  assign dataMem_6_7__T_74_addr = dataMem_6_7__T_74_addr_pipe_0;
  assign dataMem_6_7__T_74_data = dataMem_6_7[dataMem_6_7__T_74_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_7__T_178_addr = dataMem_6_7__T_178_addr_pipe_0;
  assign dataMem_6_7__T_178_data = dataMem_6_7[dataMem_6_7__T_178_addr]; // @[AXICache.scala 721:45]
  assign dataMem_6_7__T_395_data = wdata[447:440];
  assign dataMem_6_7__T_395_addr = addr_reg[13:6];
  assign dataMem_6_7__T_395_mask = wmask[55];
  assign dataMem_6_7__T_395_en = _T_100 | is_alloc;
  assign dataMem_7_0__T_84_addr = dataMem_7_0__T_84_addr_pipe_0;
  assign dataMem_7_0__T_84_data = dataMem_7_0[dataMem_7_0__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_0__T_189_addr = dataMem_7_0__T_189_addr_pipe_0;
  assign dataMem_7_0__T_189_data = dataMem_7_0[dataMem_7_0__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_0__T_414_data = wdata[455:448];
  assign dataMem_7_0__T_414_addr = addr_reg[13:6];
  assign dataMem_7_0__T_414_mask = wmask[56];
  assign dataMem_7_0__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_1__T_84_addr = dataMem_7_1__T_84_addr_pipe_0;
  assign dataMem_7_1__T_84_data = dataMem_7_1[dataMem_7_1__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_1__T_189_addr = dataMem_7_1__T_189_addr_pipe_0;
  assign dataMem_7_1__T_189_data = dataMem_7_1[dataMem_7_1__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_1__T_414_data = wdata[463:456];
  assign dataMem_7_1__T_414_addr = addr_reg[13:6];
  assign dataMem_7_1__T_414_mask = wmask[57];
  assign dataMem_7_1__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_2__T_84_addr = dataMem_7_2__T_84_addr_pipe_0;
  assign dataMem_7_2__T_84_data = dataMem_7_2[dataMem_7_2__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_2__T_189_addr = dataMem_7_2__T_189_addr_pipe_0;
  assign dataMem_7_2__T_189_data = dataMem_7_2[dataMem_7_2__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_2__T_414_data = wdata[471:464];
  assign dataMem_7_2__T_414_addr = addr_reg[13:6];
  assign dataMem_7_2__T_414_mask = wmask[58];
  assign dataMem_7_2__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_3__T_84_addr = dataMem_7_3__T_84_addr_pipe_0;
  assign dataMem_7_3__T_84_data = dataMem_7_3[dataMem_7_3__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_3__T_189_addr = dataMem_7_3__T_189_addr_pipe_0;
  assign dataMem_7_3__T_189_data = dataMem_7_3[dataMem_7_3__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_3__T_414_data = wdata[479:472];
  assign dataMem_7_3__T_414_addr = addr_reg[13:6];
  assign dataMem_7_3__T_414_mask = wmask[59];
  assign dataMem_7_3__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_4__T_84_addr = dataMem_7_4__T_84_addr_pipe_0;
  assign dataMem_7_4__T_84_data = dataMem_7_4[dataMem_7_4__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_4__T_189_addr = dataMem_7_4__T_189_addr_pipe_0;
  assign dataMem_7_4__T_189_data = dataMem_7_4[dataMem_7_4__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_4__T_414_data = wdata[487:480];
  assign dataMem_7_4__T_414_addr = addr_reg[13:6];
  assign dataMem_7_4__T_414_mask = wmask[60];
  assign dataMem_7_4__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_5__T_84_addr = dataMem_7_5__T_84_addr_pipe_0;
  assign dataMem_7_5__T_84_data = dataMem_7_5[dataMem_7_5__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_5__T_189_addr = dataMem_7_5__T_189_addr_pipe_0;
  assign dataMem_7_5__T_189_data = dataMem_7_5[dataMem_7_5__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_5__T_414_data = wdata[495:488];
  assign dataMem_7_5__T_414_addr = addr_reg[13:6];
  assign dataMem_7_5__T_414_mask = wmask[61];
  assign dataMem_7_5__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_6__T_84_addr = dataMem_7_6__T_84_addr_pipe_0;
  assign dataMem_7_6__T_84_data = dataMem_7_6[dataMem_7_6__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_6__T_189_addr = dataMem_7_6__T_189_addr_pipe_0;
  assign dataMem_7_6__T_189_data = dataMem_7_6[dataMem_7_6__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_6__T_414_data = wdata[503:496];
  assign dataMem_7_6__T_414_addr = addr_reg[13:6];
  assign dataMem_7_6__T_414_mask = wmask[62];
  assign dataMem_7_6__T_414_en = _T_100 | is_alloc;
  assign dataMem_7_7__T_84_addr = dataMem_7_7__T_84_addr_pipe_0;
  assign dataMem_7_7__T_84_data = dataMem_7_7[dataMem_7_7__T_84_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_7__T_189_addr = dataMem_7_7__T_189_addr_pipe_0;
  assign dataMem_7_7__T_189_data = dataMem_7_7[dataMem_7_7__T_189_addr]; // @[AXICache.scala 721:45]
  assign dataMem_7_7__T_414_data = wdata[511:504];
  assign dataMem_7_7__T_414_addr = addr_reg[13:6];
  assign dataMem_7_7__T_414_mask = wmask[63];
  assign dataMem_7_7__T_414_en = _T_100 | is_alloc;
  assign io_cpu_flush_done = _T_480 ? 1'h0 : _GEN_395; // @[AXICache.scala 850:21 AXICache.scala 924:27]
  assign io_cpu_req_ready = is_idle | _T_216; // @[AXICache.scala 765:20]
  assign io_cpu_resp_valid = _T_217 | _T_231; // @[AXICache.scala 769:21]
  assign io_cpu_resp_bits_data = 3'h7 == off_reg ? read[511:448] : _GEN_25; // @[AXICache.scala 768:25]
  assign io_cpu_resp_bits_tag = cpu_tag_reg; // @[AXICache.scala 771:24]
  assign io_mem_rd_cmd_valid = _T_480 ? _GEN_373 : _GEN_399; // @[AXICache.scala 814:23 AXICache.scala 869:29 AXICache.scala 882:29 AXICache.scala 902:27 AXICache.scala 956:27]
  assign io_mem_rd_cmd_bits_addr = _T_416[31:0]; // @[AXICache.scala 812:27]
  assign io_mem_rd_data_ready = state == 3'h6; // @[AXICache.scala 817:24]
  assign io_mem_wr_cmd_valid = _T_480 ? _GEN_372 : _GEN_398; // @[AXICache.scala 837:23 AXICache.scala 868:29 AXICache.scala 881:29 AXICache.scala 955:27]
  assign io_mem_wr_cmd_bits_addr = _T_434[31:0]; // @[AXICache.scala 835:27]
  assign io_mem_wr_data_valid = _T_480 ? _GEN_374 : _GEN_400; // @[AXICache.scala 847:24 AXICache.scala 891:28 AXICache.scala 966:28]
  assign io_mem_wr_data_bits = flush_mode ? _GEN_330 : _GEN_338; // @[AXICache.scala 840:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    metaMem_tag[initvar] = _RAND_0[49:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_0[initvar] = _RAND_5[7:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_1[initvar] = _RAND_9[7:0];
  _RAND_13 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_2[initvar] = _RAND_13[7:0];
  _RAND_17 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_3[initvar] = _RAND_17[7:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_4[initvar] = _RAND_21[7:0];
  _RAND_25 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_5[initvar] = _RAND_25[7:0];
  _RAND_29 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_6[initvar] = _RAND_29[7:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_0_7[initvar] = _RAND_33[7:0];
  _RAND_37 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_0[initvar] = _RAND_37[7:0];
  _RAND_41 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_1[initvar] = _RAND_41[7:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_2[initvar] = _RAND_45[7:0];
  _RAND_49 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_3[initvar] = _RAND_49[7:0];
  _RAND_53 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_4[initvar] = _RAND_53[7:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_5[initvar] = _RAND_57[7:0];
  _RAND_61 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_6[initvar] = _RAND_61[7:0];
  _RAND_65 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_1_7[initvar] = _RAND_65[7:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_0[initvar] = _RAND_69[7:0];
  _RAND_73 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_1[initvar] = _RAND_73[7:0];
  _RAND_77 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_2[initvar] = _RAND_77[7:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_3[initvar] = _RAND_81[7:0];
  _RAND_85 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_4[initvar] = _RAND_85[7:0];
  _RAND_89 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_5[initvar] = _RAND_89[7:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_6[initvar] = _RAND_93[7:0];
  _RAND_97 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_2_7[initvar] = _RAND_97[7:0];
  _RAND_101 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_0[initvar] = _RAND_101[7:0];
  _RAND_105 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_1[initvar] = _RAND_105[7:0];
  _RAND_109 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_2[initvar] = _RAND_109[7:0];
  _RAND_113 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_3[initvar] = _RAND_113[7:0];
  _RAND_117 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_4[initvar] = _RAND_117[7:0];
  _RAND_121 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_5[initvar] = _RAND_121[7:0];
  _RAND_125 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_6[initvar] = _RAND_125[7:0];
  _RAND_129 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_3_7[initvar] = _RAND_129[7:0];
  _RAND_133 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_0[initvar] = _RAND_133[7:0];
  _RAND_137 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_1[initvar] = _RAND_137[7:0];
  _RAND_141 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_2[initvar] = _RAND_141[7:0];
  _RAND_145 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_3[initvar] = _RAND_145[7:0];
  _RAND_149 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_4[initvar] = _RAND_149[7:0];
  _RAND_153 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_5[initvar] = _RAND_153[7:0];
  _RAND_157 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_6[initvar] = _RAND_157[7:0];
  _RAND_161 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_4_7[initvar] = _RAND_161[7:0];
  _RAND_165 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_0[initvar] = _RAND_165[7:0];
  _RAND_169 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_1[initvar] = _RAND_169[7:0];
  _RAND_173 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_2[initvar] = _RAND_173[7:0];
  _RAND_177 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_3[initvar] = _RAND_177[7:0];
  _RAND_181 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_4[initvar] = _RAND_181[7:0];
  _RAND_185 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_5[initvar] = _RAND_185[7:0];
  _RAND_189 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_6[initvar] = _RAND_189[7:0];
  _RAND_193 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_5_7[initvar] = _RAND_193[7:0];
  _RAND_197 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_0[initvar] = _RAND_197[7:0];
  _RAND_201 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_1[initvar] = _RAND_201[7:0];
  _RAND_205 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_2[initvar] = _RAND_205[7:0];
  _RAND_209 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_3[initvar] = _RAND_209[7:0];
  _RAND_213 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_4[initvar] = _RAND_213[7:0];
  _RAND_217 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_5[initvar] = _RAND_217[7:0];
  _RAND_221 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_6[initvar] = _RAND_221[7:0];
  _RAND_225 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_6_7[initvar] = _RAND_225[7:0];
  _RAND_229 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_0[initvar] = _RAND_229[7:0];
  _RAND_233 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_1[initvar] = _RAND_233[7:0];
  _RAND_237 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_2[initvar] = _RAND_237[7:0];
  _RAND_241 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_3[initvar] = _RAND_241[7:0];
  _RAND_245 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_4[initvar] = _RAND_245[7:0];
  _RAND_249 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_5[initvar] = _RAND_249[7:0];
  _RAND_253 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_6[initvar] = _RAND_253[7:0];
  _RAND_257 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    dataMem_7_7[initvar] = _RAND_257[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  metaMem_tag_rmeta_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  metaMem_tag_rmeta_addr_pipe_0 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  metaMem_tag__T_431_en_pipe_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  metaMem_tag__T_431_addr_pipe_0 = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  dataMem_0_0__T_14_addr_pipe_0 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  dataMem_0_0__T_112_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dataMem_0_0__T_112_addr_pipe_0 = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  dataMem_0_1__T_14_addr_pipe_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  dataMem_0_1__T_112_en_pipe_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  dataMem_0_1__T_112_addr_pipe_0 = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  dataMem_0_2__T_14_addr_pipe_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  dataMem_0_2__T_112_en_pipe_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dataMem_0_2__T_112_addr_pipe_0 = _RAND_16[7:0];
  _RAND_18 = {1{`RANDOM}};
  dataMem_0_3__T_14_addr_pipe_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  dataMem_0_3__T_112_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dataMem_0_3__T_112_addr_pipe_0 = _RAND_20[7:0];
  _RAND_22 = {1{`RANDOM}};
  dataMem_0_4__T_14_addr_pipe_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  dataMem_0_4__T_112_en_pipe_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  dataMem_0_4__T_112_addr_pipe_0 = _RAND_24[7:0];
  _RAND_26 = {1{`RANDOM}};
  dataMem_0_5__T_14_addr_pipe_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  dataMem_0_5__T_112_en_pipe_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  dataMem_0_5__T_112_addr_pipe_0 = _RAND_28[7:0];
  _RAND_30 = {1{`RANDOM}};
  dataMem_0_6__T_14_addr_pipe_0 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  dataMem_0_6__T_112_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dataMem_0_6__T_112_addr_pipe_0 = _RAND_32[7:0];
  _RAND_34 = {1{`RANDOM}};
  dataMem_0_7__T_14_addr_pipe_0 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  dataMem_0_7__T_112_en_pipe_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  dataMem_0_7__T_112_addr_pipe_0 = _RAND_36[7:0];
  _RAND_38 = {1{`RANDOM}};
  dataMem_1_0__T_24_addr_pipe_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  dataMem_1_0__T_123_en_pipe_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  dataMem_1_0__T_123_addr_pipe_0 = _RAND_40[7:0];
  _RAND_42 = {1{`RANDOM}};
  dataMem_1_1__T_24_addr_pipe_0 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  dataMem_1_1__T_123_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  dataMem_1_1__T_123_addr_pipe_0 = _RAND_44[7:0];
  _RAND_46 = {1{`RANDOM}};
  dataMem_1_2__T_24_addr_pipe_0 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  dataMem_1_2__T_123_en_pipe_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  dataMem_1_2__T_123_addr_pipe_0 = _RAND_48[7:0];
  _RAND_50 = {1{`RANDOM}};
  dataMem_1_3__T_24_addr_pipe_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  dataMem_1_3__T_123_en_pipe_0 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  dataMem_1_3__T_123_addr_pipe_0 = _RAND_52[7:0];
  _RAND_54 = {1{`RANDOM}};
  dataMem_1_4__T_24_addr_pipe_0 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  dataMem_1_4__T_123_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  dataMem_1_4__T_123_addr_pipe_0 = _RAND_56[7:0];
  _RAND_58 = {1{`RANDOM}};
  dataMem_1_5__T_24_addr_pipe_0 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  dataMem_1_5__T_123_en_pipe_0 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  dataMem_1_5__T_123_addr_pipe_0 = _RAND_60[7:0];
  _RAND_62 = {1{`RANDOM}};
  dataMem_1_6__T_24_addr_pipe_0 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  dataMem_1_6__T_123_en_pipe_0 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  dataMem_1_6__T_123_addr_pipe_0 = _RAND_64[7:0];
  _RAND_66 = {1{`RANDOM}};
  dataMem_1_7__T_24_addr_pipe_0 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  dataMem_1_7__T_123_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dataMem_1_7__T_123_addr_pipe_0 = _RAND_68[7:0];
  _RAND_70 = {1{`RANDOM}};
  dataMem_2_0__T_34_addr_pipe_0 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  dataMem_2_0__T_134_en_pipe_0 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dataMem_2_0__T_134_addr_pipe_0 = _RAND_72[7:0];
  _RAND_74 = {1{`RANDOM}};
  dataMem_2_1__T_34_addr_pipe_0 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  dataMem_2_1__T_134_en_pipe_0 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dataMem_2_1__T_134_addr_pipe_0 = _RAND_76[7:0];
  _RAND_78 = {1{`RANDOM}};
  dataMem_2_2__T_34_addr_pipe_0 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  dataMem_2_2__T_134_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dataMem_2_2__T_134_addr_pipe_0 = _RAND_80[7:0];
  _RAND_82 = {1{`RANDOM}};
  dataMem_2_3__T_34_addr_pipe_0 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  dataMem_2_3__T_134_en_pipe_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dataMem_2_3__T_134_addr_pipe_0 = _RAND_84[7:0];
  _RAND_86 = {1{`RANDOM}};
  dataMem_2_4__T_34_addr_pipe_0 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  dataMem_2_4__T_134_en_pipe_0 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dataMem_2_4__T_134_addr_pipe_0 = _RAND_88[7:0];
  _RAND_90 = {1{`RANDOM}};
  dataMem_2_5__T_34_addr_pipe_0 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  dataMem_2_5__T_134_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dataMem_2_5__T_134_addr_pipe_0 = _RAND_92[7:0];
  _RAND_94 = {1{`RANDOM}};
  dataMem_2_6__T_34_addr_pipe_0 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  dataMem_2_6__T_134_en_pipe_0 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dataMem_2_6__T_134_addr_pipe_0 = _RAND_96[7:0];
  _RAND_98 = {1{`RANDOM}};
  dataMem_2_7__T_34_addr_pipe_0 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  dataMem_2_7__T_134_en_pipe_0 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dataMem_2_7__T_134_addr_pipe_0 = _RAND_100[7:0];
  _RAND_102 = {1{`RANDOM}};
  dataMem_3_0__T_44_addr_pipe_0 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  dataMem_3_0__T_145_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dataMem_3_0__T_145_addr_pipe_0 = _RAND_104[7:0];
  _RAND_106 = {1{`RANDOM}};
  dataMem_3_1__T_44_addr_pipe_0 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  dataMem_3_1__T_145_en_pipe_0 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dataMem_3_1__T_145_addr_pipe_0 = _RAND_108[7:0];
  _RAND_110 = {1{`RANDOM}};
  dataMem_3_2__T_44_addr_pipe_0 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  dataMem_3_2__T_145_en_pipe_0 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dataMem_3_2__T_145_addr_pipe_0 = _RAND_112[7:0];
  _RAND_114 = {1{`RANDOM}};
  dataMem_3_3__T_44_addr_pipe_0 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  dataMem_3_3__T_145_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dataMem_3_3__T_145_addr_pipe_0 = _RAND_116[7:0];
  _RAND_118 = {1{`RANDOM}};
  dataMem_3_4__T_44_addr_pipe_0 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  dataMem_3_4__T_145_en_pipe_0 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dataMem_3_4__T_145_addr_pipe_0 = _RAND_120[7:0];
  _RAND_122 = {1{`RANDOM}};
  dataMem_3_5__T_44_addr_pipe_0 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  dataMem_3_5__T_145_en_pipe_0 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dataMem_3_5__T_145_addr_pipe_0 = _RAND_124[7:0];
  _RAND_126 = {1{`RANDOM}};
  dataMem_3_6__T_44_addr_pipe_0 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  dataMem_3_6__T_145_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dataMem_3_6__T_145_addr_pipe_0 = _RAND_128[7:0];
  _RAND_130 = {1{`RANDOM}};
  dataMem_3_7__T_44_addr_pipe_0 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  dataMem_3_7__T_145_en_pipe_0 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  dataMem_3_7__T_145_addr_pipe_0 = _RAND_132[7:0];
  _RAND_134 = {1{`RANDOM}};
  dataMem_4_0__T_54_addr_pipe_0 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  dataMem_4_0__T_156_en_pipe_0 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  dataMem_4_0__T_156_addr_pipe_0 = _RAND_136[7:0];
  _RAND_138 = {1{`RANDOM}};
  dataMem_4_1__T_54_addr_pipe_0 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  dataMem_4_1__T_156_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  dataMem_4_1__T_156_addr_pipe_0 = _RAND_140[7:0];
  _RAND_142 = {1{`RANDOM}};
  dataMem_4_2__T_54_addr_pipe_0 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  dataMem_4_2__T_156_en_pipe_0 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  dataMem_4_2__T_156_addr_pipe_0 = _RAND_144[7:0];
  _RAND_146 = {1{`RANDOM}};
  dataMem_4_3__T_54_addr_pipe_0 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  dataMem_4_3__T_156_en_pipe_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  dataMem_4_3__T_156_addr_pipe_0 = _RAND_148[7:0];
  _RAND_150 = {1{`RANDOM}};
  dataMem_4_4__T_54_addr_pipe_0 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  dataMem_4_4__T_156_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  dataMem_4_4__T_156_addr_pipe_0 = _RAND_152[7:0];
  _RAND_154 = {1{`RANDOM}};
  dataMem_4_5__T_54_addr_pipe_0 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  dataMem_4_5__T_156_en_pipe_0 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  dataMem_4_5__T_156_addr_pipe_0 = _RAND_156[7:0];
  _RAND_158 = {1{`RANDOM}};
  dataMem_4_6__T_54_addr_pipe_0 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  dataMem_4_6__T_156_en_pipe_0 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  dataMem_4_6__T_156_addr_pipe_0 = _RAND_160[7:0];
  _RAND_162 = {1{`RANDOM}};
  dataMem_4_7__T_54_addr_pipe_0 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  dataMem_4_7__T_156_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  dataMem_4_7__T_156_addr_pipe_0 = _RAND_164[7:0];
  _RAND_166 = {1{`RANDOM}};
  dataMem_5_0__T_64_addr_pipe_0 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  dataMem_5_0__T_167_en_pipe_0 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  dataMem_5_0__T_167_addr_pipe_0 = _RAND_168[7:0];
  _RAND_170 = {1{`RANDOM}};
  dataMem_5_1__T_64_addr_pipe_0 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  dataMem_5_1__T_167_en_pipe_0 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  dataMem_5_1__T_167_addr_pipe_0 = _RAND_172[7:0];
  _RAND_174 = {1{`RANDOM}};
  dataMem_5_2__T_64_addr_pipe_0 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  dataMem_5_2__T_167_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  dataMem_5_2__T_167_addr_pipe_0 = _RAND_176[7:0];
  _RAND_178 = {1{`RANDOM}};
  dataMem_5_3__T_64_addr_pipe_0 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  dataMem_5_3__T_167_en_pipe_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  dataMem_5_3__T_167_addr_pipe_0 = _RAND_180[7:0];
  _RAND_182 = {1{`RANDOM}};
  dataMem_5_4__T_64_addr_pipe_0 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  dataMem_5_4__T_167_en_pipe_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  dataMem_5_4__T_167_addr_pipe_0 = _RAND_184[7:0];
  _RAND_186 = {1{`RANDOM}};
  dataMem_5_5__T_64_addr_pipe_0 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  dataMem_5_5__T_167_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  dataMem_5_5__T_167_addr_pipe_0 = _RAND_188[7:0];
  _RAND_190 = {1{`RANDOM}};
  dataMem_5_6__T_64_addr_pipe_0 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  dataMem_5_6__T_167_en_pipe_0 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  dataMem_5_6__T_167_addr_pipe_0 = _RAND_192[7:0];
  _RAND_194 = {1{`RANDOM}};
  dataMem_5_7__T_64_addr_pipe_0 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  dataMem_5_7__T_167_en_pipe_0 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  dataMem_5_7__T_167_addr_pipe_0 = _RAND_196[7:0];
  _RAND_198 = {1{`RANDOM}};
  dataMem_6_0__T_74_addr_pipe_0 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  dataMem_6_0__T_178_en_pipe_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  dataMem_6_0__T_178_addr_pipe_0 = _RAND_200[7:0];
  _RAND_202 = {1{`RANDOM}};
  dataMem_6_1__T_74_addr_pipe_0 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  dataMem_6_1__T_178_en_pipe_0 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  dataMem_6_1__T_178_addr_pipe_0 = _RAND_204[7:0];
  _RAND_206 = {1{`RANDOM}};
  dataMem_6_2__T_74_addr_pipe_0 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  dataMem_6_2__T_178_en_pipe_0 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  dataMem_6_2__T_178_addr_pipe_0 = _RAND_208[7:0];
  _RAND_210 = {1{`RANDOM}};
  dataMem_6_3__T_74_addr_pipe_0 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  dataMem_6_3__T_178_en_pipe_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  dataMem_6_3__T_178_addr_pipe_0 = _RAND_212[7:0];
  _RAND_214 = {1{`RANDOM}};
  dataMem_6_4__T_74_addr_pipe_0 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  dataMem_6_4__T_178_en_pipe_0 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  dataMem_6_4__T_178_addr_pipe_0 = _RAND_216[7:0];
  _RAND_218 = {1{`RANDOM}};
  dataMem_6_5__T_74_addr_pipe_0 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  dataMem_6_5__T_178_en_pipe_0 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  dataMem_6_5__T_178_addr_pipe_0 = _RAND_220[7:0];
  _RAND_222 = {1{`RANDOM}};
  dataMem_6_6__T_74_addr_pipe_0 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  dataMem_6_6__T_178_en_pipe_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  dataMem_6_6__T_178_addr_pipe_0 = _RAND_224[7:0];
  _RAND_226 = {1{`RANDOM}};
  dataMem_6_7__T_74_addr_pipe_0 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  dataMem_6_7__T_178_en_pipe_0 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  dataMem_6_7__T_178_addr_pipe_0 = _RAND_228[7:0];
  _RAND_230 = {1{`RANDOM}};
  dataMem_7_0__T_84_addr_pipe_0 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  dataMem_7_0__T_189_en_pipe_0 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  dataMem_7_0__T_189_addr_pipe_0 = _RAND_232[7:0];
  _RAND_234 = {1{`RANDOM}};
  dataMem_7_1__T_84_addr_pipe_0 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  dataMem_7_1__T_189_en_pipe_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  dataMem_7_1__T_189_addr_pipe_0 = _RAND_236[7:0];
  _RAND_238 = {1{`RANDOM}};
  dataMem_7_2__T_84_addr_pipe_0 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  dataMem_7_2__T_189_en_pipe_0 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  dataMem_7_2__T_189_addr_pipe_0 = _RAND_240[7:0];
  _RAND_242 = {1{`RANDOM}};
  dataMem_7_3__T_84_addr_pipe_0 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  dataMem_7_3__T_189_en_pipe_0 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  dataMem_7_3__T_189_addr_pipe_0 = _RAND_244[7:0];
  _RAND_246 = {1{`RANDOM}};
  dataMem_7_4__T_84_addr_pipe_0 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  dataMem_7_4__T_189_en_pipe_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  dataMem_7_4__T_189_addr_pipe_0 = _RAND_248[7:0];
  _RAND_250 = {1{`RANDOM}};
  dataMem_7_5__T_84_addr_pipe_0 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  dataMem_7_5__T_189_en_pipe_0 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  dataMem_7_5__T_189_addr_pipe_0 = _RAND_252[7:0];
  _RAND_254 = {1{`RANDOM}};
  dataMem_7_6__T_84_addr_pipe_0 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  dataMem_7_6__T_189_en_pipe_0 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  dataMem_7_6__T_189_addr_pipe_0 = _RAND_256[7:0];
  _RAND_258 = {1{`RANDOM}};
  dataMem_7_7__T_84_addr_pipe_0 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  dataMem_7_7__T_189_en_pipe_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  dataMem_7_7__T_189_addr_pipe_0 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  state = _RAND_261[2:0];
  _RAND_262 = {1{`RANDOM}};
  flush_state = _RAND_262[2:0];
  _RAND_263 = {1{`RANDOM}};
  flush_mode = _RAND_263[0:0];
  _RAND_264 = {8{`RANDOM}};
  v = _RAND_264[255:0];
  _RAND_265 = {8{`RANDOM}};
  d = _RAND_265[255:0];
  _RAND_266 = {2{`RANDOM}};
  addr_reg = _RAND_266[63:0];
  _RAND_267 = {1{`RANDOM}};
  cpu_tag_reg = _RAND_267[7:0];
  _RAND_268 = {2{`RANDOM}};
  cpu_data = _RAND_268[63:0];
  _RAND_269 = {1{`RANDOM}};
  cpu_mask = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  read_count = _RAND_270[2:0];
  _RAND_271 = {1{`RANDOM}};
  write_count = _RAND_271[2:0];
  _RAND_272 = {1{`RANDOM}};
  set_count = _RAND_272[7:0];
  _RAND_273 = {2{`RANDOM}};
  block_rmeta_tag = _RAND_273[49:0];
  _RAND_274 = {1{`RANDOM}};
  is_alloc_reg = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ren_reg = _RAND_275[0:0];
  _RAND_276 = {16{`RANDOM}};
  rdata_buf = _RAND_276[511:0];
  _RAND_277 = {2{`RANDOM}};
  refill_buf_0 = _RAND_277[63:0];
  _RAND_278 = {2{`RANDOM}};
  refill_buf_1 = _RAND_278[63:0];
  _RAND_279 = {2{`RANDOM}};
  refill_buf_2 = _RAND_279[63:0];
  _RAND_280 = {2{`RANDOM}};
  refill_buf_3 = _RAND_280[63:0];
  _RAND_281 = {2{`RANDOM}};
  refill_buf_4 = _RAND_281[63:0];
  _RAND_282 = {2{`RANDOM}};
  refill_buf_5 = _RAND_282[63:0];
  _RAND_283 = {2{`RANDOM}};
  refill_buf_6 = _RAND_283[63:0];
  _RAND_284 = {2{`RANDOM}};
  refill_buf_7 = _RAND_284[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(metaMem_tag__T_262_en & metaMem_tag__T_262_mask) begin
      metaMem_tag[metaMem_tag__T_262_addr] <= metaMem_tag__T_262_data; // @[AXICache.scala 720:28]
    end
    metaMem_tag_rmeta_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      metaMem_tag_rmeta_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    metaMem_tag__T_431_en_pipe_0 <= is_block_dirty & _T_8;
    if (is_block_dirty & _T_8) begin
      metaMem_tag__T_431_addr_pipe_0 <= set_count;
    end
    if(dataMem_0_0__T_281_en & dataMem_0_0__T_281_mask) begin
      dataMem_0_0[dataMem_0_0__T_281_addr] <= dataMem_0_0__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_0__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_0__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_0__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_1__T_281_en & dataMem_0_1__T_281_mask) begin
      dataMem_0_1[dataMem_0_1__T_281_addr] <= dataMem_0_1__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_1__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_1__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_1__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_2__T_281_en & dataMem_0_2__T_281_mask) begin
      dataMem_0_2[dataMem_0_2__T_281_addr] <= dataMem_0_2__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_2__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_2__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_2__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_3__T_281_en & dataMem_0_3__T_281_mask) begin
      dataMem_0_3[dataMem_0_3__T_281_addr] <= dataMem_0_3__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_3__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_3__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_3__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_4__T_281_en & dataMem_0_4__T_281_mask) begin
      dataMem_0_4[dataMem_0_4__T_281_addr] <= dataMem_0_4__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_4__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_4__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_4__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_5__T_281_en & dataMem_0_5__T_281_mask) begin
      dataMem_0_5[dataMem_0_5__T_281_addr] <= dataMem_0_5__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_5__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_5__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_5__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_6__T_281_en & dataMem_0_6__T_281_mask) begin
      dataMem_0_6[dataMem_0_6__T_281_addr] <= dataMem_0_6__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_6__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_6__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_6__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_0_7__T_281_en & dataMem_0_7__T_281_mask) begin
      dataMem_0_7[dataMem_0_7__T_281_addr] <= dataMem_0_7__T_281_data; // @[AXICache.scala 721:45]
    end
    dataMem_0_7__T_14_addr_pipe_0 <= set_count - 8'h1;
    dataMem_0_7__T_112_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_0_7__T_112_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_0__T_300_en & dataMem_1_0__T_300_mask) begin
      dataMem_1_0[dataMem_1_0__T_300_addr] <= dataMem_1_0__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_0__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_0__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_0__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_1__T_300_en & dataMem_1_1__T_300_mask) begin
      dataMem_1_1[dataMem_1_1__T_300_addr] <= dataMem_1_1__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_1__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_1__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_1__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_2__T_300_en & dataMem_1_2__T_300_mask) begin
      dataMem_1_2[dataMem_1_2__T_300_addr] <= dataMem_1_2__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_2__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_2__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_2__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_3__T_300_en & dataMem_1_3__T_300_mask) begin
      dataMem_1_3[dataMem_1_3__T_300_addr] <= dataMem_1_3__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_3__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_3__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_3__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_4__T_300_en & dataMem_1_4__T_300_mask) begin
      dataMem_1_4[dataMem_1_4__T_300_addr] <= dataMem_1_4__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_4__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_4__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_4__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_5__T_300_en & dataMem_1_5__T_300_mask) begin
      dataMem_1_5[dataMem_1_5__T_300_addr] <= dataMem_1_5__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_5__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_5__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_5__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_6__T_300_en & dataMem_1_6__T_300_mask) begin
      dataMem_1_6[dataMem_1_6__T_300_addr] <= dataMem_1_6__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_6__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_6__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_6__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_1_7__T_300_en & dataMem_1_7__T_300_mask) begin
      dataMem_1_7[dataMem_1_7__T_300_addr] <= dataMem_1_7__T_300_data; // @[AXICache.scala 721:45]
    end
    dataMem_1_7__T_24_addr_pipe_0 <= set_count - 8'h1;
    dataMem_1_7__T_123_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_1_7__T_123_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_0__T_319_en & dataMem_2_0__T_319_mask) begin
      dataMem_2_0[dataMem_2_0__T_319_addr] <= dataMem_2_0__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_0__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_0__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_0__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_1__T_319_en & dataMem_2_1__T_319_mask) begin
      dataMem_2_1[dataMem_2_1__T_319_addr] <= dataMem_2_1__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_1__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_1__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_1__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_2__T_319_en & dataMem_2_2__T_319_mask) begin
      dataMem_2_2[dataMem_2_2__T_319_addr] <= dataMem_2_2__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_2__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_2__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_2__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_3__T_319_en & dataMem_2_3__T_319_mask) begin
      dataMem_2_3[dataMem_2_3__T_319_addr] <= dataMem_2_3__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_3__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_3__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_3__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_4__T_319_en & dataMem_2_4__T_319_mask) begin
      dataMem_2_4[dataMem_2_4__T_319_addr] <= dataMem_2_4__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_4__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_4__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_4__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_5__T_319_en & dataMem_2_5__T_319_mask) begin
      dataMem_2_5[dataMem_2_5__T_319_addr] <= dataMem_2_5__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_5__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_5__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_5__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_6__T_319_en & dataMem_2_6__T_319_mask) begin
      dataMem_2_6[dataMem_2_6__T_319_addr] <= dataMem_2_6__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_6__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_6__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_6__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_2_7__T_319_en & dataMem_2_7__T_319_mask) begin
      dataMem_2_7[dataMem_2_7__T_319_addr] <= dataMem_2_7__T_319_data; // @[AXICache.scala 721:45]
    end
    dataMem_2_7__T_34_addr_pipe_0 <= set_count - 8'h1;
    dataMem_2_7__T_134_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_2_7__T_134_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_0__T_338_en & dataMem_3_0__T_338_mask) begin
      dataMem_3_0[dataMem_3_0__T_338_addr] <= dataMem_3_0__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_0__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_0__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_0__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_1__T_338_en & dataMem_3_1__T_338_mask) begin
      dataMem_3_1[dataMem_3_1__T_338_addr] <= dataMem_3_1__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_1__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_1__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_1__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_2__T_338_en & dataMem_3_2__T_338_mask) begin
      dataMem_3_2[dataMem_3_2__T_338_addr] <= dataMem_3_2__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_2__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_2__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_2__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_3__T_338_en & dataMem_3_3__T_338_mask) begin
      dataMem_3_3[dataMem_3_3__T_338_addr] <= dataMem_3_3__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_3__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_3__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_3__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_4__T_338_en & dataMem_3_4__T_338_mask) begin
      dataMem_3_4[dataMem_3_4__T_338_addr] <= dataMem_3_4__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_4__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_4__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_4__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_5__T_338_en & dataMem_3_5__T_338_mask) begin
      dataMem_3_5[dataMem_3_5__T_338_addr] <= dataMem_3_5__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_5__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_5__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_5__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_6__T_338_en & dataMem_3_6__T_338_mask) begin
      dataMem_3_6[dataMem_3_6__T_338_addr] <= dataMem_3_6__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_6__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_6__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_6__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_3_7__T_338_en & dataMem_3_7__T_338_mask) begin
      dataMem_3_7[dataMem_3_7__T_338_addr] <= dataMem_3_7__T_338_data; // @[AXICache.scala 721:45]
    end
    dataMem_3_7__T_44_addr_pipe_0 <= set_count - 8'h1;
    dataMem_3_7__T_145_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_3_7__T_145_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_0__T_357_en & dataMem_4_0__T_357_mask) begin
      dataMem_4_0[dataMem_4_0__T_357_addr] <= dataMem_4_0__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_0__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_0__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_0__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_1__T_357_en & dataMem_4_1__T_357_mask) begin
      dataMem_4_1[dataMem_4_1__T_357_addr] <= dataMem_4_1__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_1__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_1__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_1__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_2__T_357_en & dataMem_4_2__T_357_mask) begin
      dataMem_4_2[dataMem_4_2__T_357_addr] <= dataMem_4_2__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_2__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_2__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_2__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_3__T_357_en & dataMem_4_3__T_357_mask) begin
      dataMem_4_3[dataMem_4_3__T_357_addr] <= dataMem_4_3__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_3__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_3__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_3__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_4__T_357_en & dataMem_4_4__T_357_mask) begin
      dataMem_4_4[dataMem_4_4__T_357_addr] <= dataMem_4_4__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_4__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_4__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_4__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_5__T_357_en & dataMem_4_5__T_357_mask) begin
      dataMem_4_5[dataMem_4_5__T_357_addr] <= dataMem_4_5__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_5__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_5__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_5__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_6__T_357_en & dataMem_4_6__T_357_mask) begin
      dataMem_4_6[dataMem_4_6__T_357_addr] <= dataMem_4_6__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_6__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_6__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_6__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_4_7__T_357_en & dataMem_4_7__T_357_mask) begin
      dataMem_4_7[dataMem_4_7__T_357_addr] <= dataMem_4_7__T_357_data; // @[AXICache.scala 721:45]
    end
    dataMem_4_7__T_54_addr_pipe_0 <= set_count - 8'h1;
    dataMem_4_7__T_156_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_4_7__T_156_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_0__T_376_en & dataMem_5_0__T_376_mask) begin
      dataMem_5_0[dataMem_5_0__T_376_addr] <= dataMem_5_0__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_0__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_0__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_0__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_1__T_376_en & dataMem_5_1__T_376_mask) begin
      dataMem_5_1[dataMem_5_1__T_376_addr] <= dataMem_5_1__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_1__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_1__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_1__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_2__T_376_en & dataMem_5_2__T_376_mask) begin
      dataMem_5_2[dataMem_5_2__T_376_addr] <= dataMem_5_2__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_2__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_2__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_2__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_3__T_376_en & dataMem_5_3__T_376_mask) begin
      dataMem_5_3[dataMem_5_3__T_376_addr] <= dataMem_5_3__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_3__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_3__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_3__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_4__T_376_en & dataMem_5_4__T_376_mask) begin
      dataMem_5_4[dataMem_5_4__T_376_addr] <= dataMem_5_4__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_4__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_4__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_4__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_5__T_376_en & dataMem_5_5__T_376_mask) begin
      dataMem_5_5[dataMem_5_5__T_376_addr] <= dataMem_5_5__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_5__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_5__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_5__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_6__T_376_en & dataMem_5_6__T_376_mask) begin
      dataMem_5_6[dataMem_5_6__T_376_addr] <= dataMem_5_6__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_6__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_6__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_6__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_5_7__T_376_en & dataMem_5_7__T_376_mask) begin
      dataMem_5_7[dataMem_5_7__T_376_addr] <= dataMem_5_7__T_376_data; // @[AXICache.scala 721:45]
    end
    dataMem_5_7__T_64_addr_pipe_0 <= set_count - 8'h1;
    dataMem_5_7__T_167_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_5_7__T_167_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_0__T_395_en & dataMem_6_0__T_395_mask) begin
      dataMem_6_0[dataMem_6_0__T_395_addr] <= dataMem_6_0__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_0__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_0__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_0__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_1__T_395_en & dataMem_6_1__T_395_mask) begin
      dataMem_6_1[dataMem_6_1__T_395_addr] <= dataMem_6_1__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_1__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_1__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_1__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_2__T_395_en & dataMem_6_2__T_395_mask) begin
      dataMem_6_2[dataMem_6_2__T_395_addr] <= dataMem_6_2__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_2__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_2__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_2__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_3__T_395_en & dataMem_6_3__T_395_mask) begin
      dataMem_6_3[dataMem_6_3__T_395_addr] <= dataMem_6_3__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_3__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_3__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_3__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_4__T_395_en & dataMem_6_4__T_395_mask) begin
      dataMem_6_4[dataMem_6_4__T_395_addr] <= dataMem_6_4__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_4__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_4__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_4__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_5__T_395_en & dataMem_6_5__T_395_mask) begin
      dataMem_6_5[dataMem_6_5__T_395_addr] <= dataMem_6_5__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_5__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_5__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_5__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_6__T_395_en & dataMem_6_6__T_395_mask) begin
      dataMem_6_6[dataMem_6_6__T_395_addr] <= dataMem_6_6__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_6__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_6__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_6__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_6_7__T_395_en & dataMem_6_7__T_395_mask) begin
      dataMem_6_7[dataMem_6_7__T_395_addr] <= dataMem_6_7__T_395_data; // @[AXICache.scala 721:45]
    end
    dataMem_6_7__T_74_addr_pipe_0 <= set_count - 8'h1;
    dataMem_6_7__T_178_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_6_7__T_178_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_0__T_414_en & dataMem_7_0__T_414_mask) begin
      dataMem_7_0[dataMem_7_0__T_414_addr] <= dataMem_7_0__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_0__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_0__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_0__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_1__T_414_en & dataMem_7_1__T_414_mask) begin
      dataMem_7_1[dataMem_7_1__T_414_addr] <= dataMem_7_1__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_1__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_1__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_1__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_2__T_414_en & dataMem_7_2__T_414_mask) begin
      dataMem_7_2[dataMem_7_2__T_414_addr] <= dataMem_7_2__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_2__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_2__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_2__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_3__T_414_en & dataMem_7_3__T_414_mask) begin
      dataMem_7_3[dataMem_7_3__T_414_addr] <= dataMem_7_3__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_3__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_3__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_3__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_4__T_414_en & dataMem_7_4__T_414_mask) begin
      dataMem_7_4[dataMem_7_4__T_414_addr] <= dataMem_7_4__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_4__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_4__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_4__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_5__T_414_en & dataMem_7_5__T_414_mask) begin
      dataMem_7_5[dataMem_7_5__T_414_addr] <= dataMem_7_5__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_5__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_5__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_5__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_6__T_414_en & dataMem_7_6__T_414_mask) begin
      dataMem_7_6[dataMem_7_6__T_414_addr] <= dataMem_7_6__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_6__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_6__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_6__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if(dataMem_7_7__T_414_en & dataMem_7_7__T_414_mask) begin
      dataMem_7_7[dataMem_7_7__T_414_addr] <= dataMem_7_7__T_414_data; // @[AXICache.scala 721:45]
    end
    dataMem_7_7__T_84_addr_pipe_0 <= set_count - 8'h1;
    dataMem_7_7__T_189_en_pipe_0 <= _T_105 & io_cpu_req_valid;
    if (_T_105 & io_cpu_req_valid) begin
      dataMem_7_7__T_189_addr_pipe_0 <= io_cpu_req_bits_addr[13:6];
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_458) begin
      if (io_cpu_req_valid) begin
        if (_T_459) begin
          state <= 3'h2;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (_T_461) begin
      if (hit) begin
        if (io_cpu_req_valid) begin
          if (_T_459) begin
            state <= 3'h2;
          end else begin
            state <= 3'h1;
          end
        end else begin
          state <= 3'h0;
        end
      end else if (_T_465) begin
        state <= 3'h3;
      end else if (_T_466) begin
        state <= 3'h6;
      end
    end else if (_T_467) begin
      if (_T_99) begin
        state <= 3'h0;
      end else if (_T_465) begin
        state <= 3'h3;
      end else if (_T_466) begin
        state <= 3'h6;
      end
    end else if (_T_473) begin
      if (write_wrap_out) begin
        state <= 3'h4;
      end
    end else if (_T_474) begin
      if (io_mem_wr_ack) begin
        state <= 3'h5;
      end
    end else if (_T_475) begin
      if (_T_466) begin
        state <= 3'h6;
      end
    end else if (_T_477) begin
      if (read_wrap_out) begin
        if (_T_229) begin
          state <= 3'h2;
        end else begin
          state <= 3'h0;
        end
      end
    end
    if (reset) begin
      flush_state <= 3'h0;
    end else if (_T_480) begin
      if (io_cpu_flush) begin
        flush_state <= 3'h1;
      end
    end else if (_T_481) begin
      if (set_wrap) begin
        flush_state <= 3'h0;
      end else if (is_block_dirty) begin
        flush_state <= 3'h2;
      end
    end else if (_T_482) begin
      flush_state <= 3'h3;
    end else if (_T_483) begin
      if (_T_465) begin
        flush_state <= 3'h4;
      end
    end else if (_T_485) begin
      if (write_wrap_out) begin
        flush_state <= 3'h5;
      end
    end else if (_T_486) begin
      if (io_mem_wr_ack) begin
        flush_state <= 3'h1;
      end
    end
    if (reset) begin
      flush_mode <= 1'h0;
    end else if (_T_480) begin
      flush_mode <= _GEN_376;
    end else if (_T_481) begin
      if (set_wrap) begin
        flush_mode <= 1'h0;
      end
    end
    if (reset) begin
      v <= 256'h0;
    end else if (wen) begin
      v <= _T_250;
    end
    if (reset) begin
      d <= 256'h0;
    end else if (wen) begin
      if (_T_234) begin
        d <= _T_257;
      end else begin
        d <= _T_260;
      end
    end
    if (io_cpu_resp_valid) begin
      addr_reg <= io_cpu_req_bits_addr;
    end
    if (_T_233) begin
      cpu_tag_reg <= io_cpu_req_bits_tag;
    end
    if (io_cpu_resp_valid) begin
      cpu_data <= io_cpu_req_bits_data;
    end
    if (io_cpu_resp_valid) begin
      cpu_mask <= io_cpu_req_bits_mask;
    end
    if (reset) begin
      read_count <= 3'h0;
    end else if (_T) begin
      read_count <= _T_3;
    end
    if (reset) begin
      write_count <= 3'h0;
    end else if (_T_4) begin
      write_count <= _T_7;
    end
    if (reset) begin
      set_count <= 8'h0;
    end else if (_T_8) begin
      set_count <= _T_11;
    end
    block_rmeta_tag <= metaMem_tag__T_431_data;
    is_alloc_reg <= _T_98 & read_wrap_out;
    ren_reg <= _T_105 & io_cpu_req_valid;
    if (ren_reg) begin
      rdata_buf <= rdata;
    end
    if (_T) begin
      if (3'h0 == read_count) begin
        refill_buf_0 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h1 == read_count) begin
        refill_buf_1 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h2 == read_count) begin
        refill_buf_2 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h3 == read_count) begin
        refill_buf_3 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h4 == read_count) begin
        refill_buf_4 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h5 == read_count) begin
        refill_buf_5 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h6 == read_count) begin
        refill_buf_6 <= io_mem_rd_data_bits;
      end
    end
    if (_T) begin
      if (3'h7 == read_count) begin
        refill_buf_7 <= io_mem_rd_data_bits;
      end
    end
  end
endmodule
module Arbiter_2(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_addr,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [63:0] io_in_1_bits_addr,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [63:0] io_in_2_bits_addr,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [63:0] io_in_3_bits_addr,
  input  [63:0] io_in_3_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [63:0] io_out_bits_data,
  output [7:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [1:0]  io_chosen
);
  wire [1:0] _GEN_0 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_3 = io_in_2_valid ? 8'h2 : 8'h3; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_4 = io_in_2_valid ? 8'h0 : 8'hff; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_5 = io_in_2_valid ? 64'h0 : io_in_3_bits_data; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_6 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27]
  wire [1:0] _GEN_7 = io_in_1_valid ? 2'h1 : _GEN_0; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_10 = io_in_1_valid ? 8'h1 : _GEN_3; // @[Arbiter.scala 126:27]
  wire [7:0] _GEN_11 = io_in_1_valid ? 8'h0 : _GEN_4; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_12 = io_in_1_valid ? 64'h0 : _GEN_5; // @[Arbiter.scala 126:27]
  wire [63:0] _GEN_13 = io_in_1_valid ? io_in_1_bits_addr : _GEN_6; // @[Arbiter.scala 126:27]
  wire  _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_1 = _T | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  grant_2 = ~_T; // @[Arbiter.scala 31:78]
  wire  grant_3 = ~_T_1; // @[Arbiter.scala 31:78]
  wire  _T_6 = ~grant_3; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_2_ready = grant_2 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_3_ready = grant_3 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_6 | io_in_3_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_13; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? 64'h0 : _GEN_12; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_mask = io_in_0_valid ? 8'h0 : _GEN_11; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_out_bits_tag = io_in_0_valid ? 8'h0 : _GEN_10; // @[Arbiter.scala 124:15 Arbiter.scala 128:19 Arbiter.scala 128:19 Arbiter.scala 128:19]
  assign io_chosen = io_in_0_valid ? 2'h0 : _GEN_7; // @[Arbiter.scala 123:13 Arbiter.scala 127:17 Arbiter.scala 127:17 Arbiter.scala 127:17]
endmodule
module CacheMemoryEngine(
  input         clock,
  input         reset,
  output        io_rd_mem_0_MemReq_ready,
  input         io_rd_mem_0_MemReq_valid,
  input  [63:0] io_rd_mem_0_MemReq_bits_addr,
  output        io_rd_mem_0_MemResp_valid,
  output [63:0] io_rd_mem_0_MemResp_bits_data,
  output        io_rd_mem_1_MemReq_ready,
  input         io_rd_mem_1_MemReq_valid,
  input  [63:0] io_rd_mem_1_MemReq_bits_addr,
  output        io_rd_mem_1_MemResp_valid,
  output [63:0] io_rd_mem_1_MemResp_bits_data,
  output        io_rd_mem_2_MemReq_ready,
  input         io_rd_mem_2_MemReq_valid,
  input  [63:0] io_rd_mem_2_MemReq_bits_addr,
  output        io_rd_mem_2_MemResp_valid,
  output [63:0] io_rd_mem_2_MemResp_bits_data,
  output        io_wr_mem_0_MemReq_ready,
  input         io_wr_mem_0_MemReq_valid,
  input  [63:0] io_wr_mem_0_MemReq_bits_addr,
  input  [63:0] io_wr_mem_0_MemReq_bits_data,
  output        io_wr_mem_0_MemResp_valid,
  input         io_cache_MemReq_ready,
  output        io_cache_MemReq_valid,
  output [63:0] io_cache_MemReq_bits_addr,
  output [63:0] io_cache_MemReq_bits_data,
  output [7:0]  io_cache_MemReq_bits_mask,
  output [7:0]  io_cache_MemReq_bits_tag,
  input         io_cache_MemResp_valid,
  input  [63:0] io_cache_MemResp_bits_data,
  input  [7:0]  io_cache_MemResp_bits_tag
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  in_arb_io_in_0_ready; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_0_valid; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_in_0_bits_addr; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_1_ready; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_1_valid; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_in_1_bits_addr; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_2_ready; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_2_valid; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_in_2_bits_addr; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_3_ready; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_in_3_valid; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_in_3_bits_addr; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_in_3_bits_data; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_out_ready; // @[CacheMemoryEngine.scala 79:22]
  wire  in_arb_io_out_valid; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_out_bits_addr; // @[CacheMemoryEngine.scala 79:22]
  wire [63:0] in_arb_io_out_bits_data; // @[CacheMemoryEngine.scala 79:22]
  wire [7:0] in_arb_io_out_bits_mask; // @[CacheMemoryEngine.scala 79:22]
  wire [7:0] in_arb_io_out_bits_tag; // @[CacheMemoryEngine.scala 79:22]
  wire [1:0] in_arb_io_chosen; // @[CacheMemoryEngine.scala 79:22]
  wire  _T = in_arb_io_out_ready & in_arb_io_out_valid; // @[Decoupled.scala 40:37]
  reg [1:0] in_arb_chosen; // @[Reg.scala 15:16]
  reg [1:0] mstate; // @[CacheMemoryEngine.scala 91:23]
  wire  _T_1 = 2'h0 == mstate; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h1 == mstate; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h2 == mstate; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_13 = {{6'd0}, in_arb_chosen}; // @[CacheMemoryEngine.scala 105:52]
  wire  _T_4 = _GEN_13 == io_cache_MemResp_bits_tag; // @[CacheMemoryEngine.scala 105:52]
  wire  _T_5 = io_cache_MemResp_valid & _T_4; // @[CacheMemoryEngine.scala 105:35]
  wire  _T_6 = in_arb_chosen == 2'h0; // @[CacheMemoryEngine.scala 112:50]
  wire  _T_8 = _T_6 & _T_4; // @[CacheMemoryEngine.scala 112:59]
  wire  _T_9 = _T_8 & io_cache_MemResp_valid; // @[CacheMemoryEngine.scala 113:53]
  wire  _T_10 = mstate == 2'h2; // @[CacheMemoryEngine.scala 115:15]
  wire  _T_12 = in_arb_chosen == 2'h1; // @[CacheMemoryEngine.scala 112:50]
  wire  _T_14 = _T_12 & _T_4; // @[CacheMemoryEngine.scala 112:59]
  wire  _T_15 = _T_14 & io_cache_MemResp_valid; // @[CacheMemoryEngine.scala 113:53]
  wire  _T_18 = in_arb_chosen == 2'h2; // @[CacheMemoryEngine.scala 112:50]
  wire  _T_20 = _T_18 & _T_4; // @[CacheMemoryEngine.scala 112:59]
  wire  _T_21 = _T_20 & io_cache_MemResp_valid; // @[CacheMemoryEngine.scala 113:53]
  wire  _T_24 = in_arb_chosen == 2'h3; // @[CacheMemoryEngine.scala 120:60]
  wire  _T_26 = _T_24 & _T_4; // @[CacheMemoryEngine.scala 120:69]
  wire  _T_27 = _T_26 & io_cache_MemResp_valid; // @[CacheMemoryEngine.scala 121:53]
  reg [63:0] in_data_reg_addr; // @[Reg.scala 27:20]
  reg [63:0] in_data_reg_data; // @[Reg.scala 27:20]
  reg [7:0] in_data_reg_mask; // @[Reg.scala 27:20]
  reg [7:0] in_data_reg_tag; // @[Reg.scala 27:20]
  Arbiter_2 in_arb ( // @[CacheMemoryEngine.scala 79:22]
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_addr(in_arb_io_in_0_bits_addr),
    .io_in_1_ready(in_arb_io_in_1_ready),
    .io_in_1_valid(in_arb_io_in_1_valid),
    .io_in_1_bits_addr(in_arb_io_in_1_bits_addr),
    .io_in_2_ready(in_arb_io_in_2_ready),
    .io_in_2_valid(in_arb_io_in_2_valid),
    .io_in_2_bits_addr(in_arb_io_in_2_bits_addr),
    .io_in_3_ready(in_arb_io_in_3_ready),
    .io_in_3_valid(in_arb_io_in_3_valid),
    .io_in_3_bits_addr(in_arb_io_in_3_bits_addr),
    .io_in_3_bits_data(in_arb_io_in_3_bits_data),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_addr(in_arb_io_out_bits_addr),
    .io_out_bits_data(in_arb_io_out_bits_data),
    .io_out_bits_mask(in_arb_io_out_bits_mask),
    .io_out_bits_tag(in_arb_io_out_bits_tag),
    .io_chosen(in_arb_io_chosen)
  );
  assign io_rd_mem_0_MemReq_ready = in_arb_io_in_0_ready; // @[CacheMemoryEngine.scala 83:21]
  assign io_rd_mem_0_MemResp_valid = _T_9 & _T_10; // @[CacheMemoryEngine.scala 112:32]
  assign io_rd_mem_0_MemResp_bits_data = io_cache_MemResp_bits_data; // @[CacheMemoryEngine.scala 116:31]
  assign io_rd_mem_1_MemReq_ready = in_arb_io_in_1_ready; // @[CacheMemoryEngine.scala 83:21]
  assign io_rd_mem_1_MemResp_valid = _T_15 & _T_10; // @[CacheMemoryEngine.scala 112:32]
  assign io_rd_mem_1_MemResp_bits_data = io_cache_MemResp_bits_data; // @[CacheMemoryEngine.scala 116:31]
  assign io_rd_mem_2_MemReq_ready = in_arb_io_in_2_ready; // @[CacheMemoryEngine.scala 83:21]
  assign io_rd_mem_2_MemResp_valid = _T_21 & _T_10; // @[CacheMemoryEngine.scala 112:32]
  assign io_rd_mem_2_MemResp_bits_data = io_cache_MemResp_bits_data; // @[CacheMemoryEngine.scala 116:31]
  assign io_wr_mem_0_MemReq_ready = in_arb_io_in_3_ready; // @[CacheMemoryEngine.scala 87:31]
  assign io_wr_mem_0_MemResp_valid = _T_27 & _T_10; // @[CacheMemoryEngine.scala 120:42]
  assign io_cache_MemReq_valid = mstate == 2'h1; // @[CacheMemoryEngine.scala 130:25]
  assign io_cache_MemReq_bits_addr = in_data_reg_addr; // @[CacheMemoryEngine.scala 131:24]
  assign io_cache_MemReq_bits_data = in_data_reg_data; // @[CacheMemoryEngine.scala 131:24]
  assign io_cache_MemReq_bits_mask = in_data_reg_mask; // @[CacheMemoryEngine.scala 131:24]
  assign io_cache_MemReq_bits_tag = in_data_reg_tag; // @[CacheMemoryEngine.scala 131:24]
  assign in_arb_io_in_0_valid = io_rd_mem_0_MemReq_valid; // @[CacheMemoryEngine.scala 83:21]
  assign in_arb_io_in_0_bits_addr = io_rd_mem_0_MemReq_bits_addr; // @[CacheMemoryEngine.scala 83:21]
  assign in_arb_io_in_1_valid = io_rd_mem_1_MemReq_valid; // @[CacheMemoryEngine.scala 83:21]
  assign in_arb_io_in_1_bits_addr = io_rd_mem_1_MemReq_bits_addr; // @[CacheMemoryEngine.scala 83:21]
  assign in_arb_io_in_2_valid = io_rd_mem_2_MemReq_valid; // @[CacheMemoryEngine.scala 83:21]
  assign in_arb_io_in_2_bits_addr = io_rd_mem_2_MemReq_bits_addr; // @[CacheMemoryEngine.scala 83:21]
  assign in_arb_io_in_3_valid = io_wr_mem_0_MemReq_valid; // @[CacheMemoryEngine.scala 87:31]
  assign in_arb_io_in_3_bits_addr = io_wr_mem_0_MemReq_bits_addr; // @[CacheMemoryEngine.scala 87:31]
  assign in_arb_io_in_3_bits_data = io_wr_mem_0_MemReq_bits_data; // @[CacheMemoryEngine.scala 87:31]
  assign in_arb_io_out_ready = mstate == 2'h0; // @[CacheMemoryEngine.scala 129:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_arb_chosen = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  mstate = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  in_data_reg_addr = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  in_data_reg_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  in_data_reg_mask = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  in_data_reg_tag = _RAND_5[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (_T) begin
      in_arb_chosen <= in_arb_io_chosen;
    end
    if (reset) begin
      mstate <= 2'h0;
    end else if (_T_1) begin
      if (in_arb_io_out_valid) begin
        mstate <= 2'h1;
      end
    end else if (_T_2) begin
      if (io_cache_MemReq_ready) begin
        mstate <= 2'h2;
      end
    end else if (_T_3) begin
      if (_T_5) begin
        mstate <= 2'h0;
      end
    end
    if (reset) begin
      in_data_reg_addr <= 64'h0;
    end else if (_T) begin
      in_data_reg_addr <= in_arb_io_out_bits_addr;
    end
    if (reset) begin
      in_data_reg_data <= 64'h0;
    end else if (_T) begin
      in_data_reg_data <= in_arb_io_out_bits_data;
    end
    if (reset) begin
      in_data_reg_mask <= 8'h0;
    end else if (_T) begin
      in_data_reg_mask <= in_arb_io_out_bits_mask;
    end
    if (reset) begin
      in_data_reg_tag <= 8'h0;
    end else if (_T) begin
      in_data_reg_tag <= in_arb_io_out_bits_tag;
    end
  end
endmodule
module SplitCallDCR(
  input         clock,
  input         reset,
  output        io_In_ready,
  input         io_In_valid,
  input  [63:0] io_In_bits_dataPtrs_field2_data,
  input  [63:0] io_In_bits_dataPtrs_field1_data,
  input  [63:0] io_In_bits_dataPtrs_field0_data,
  input         io_Out_enable_ready,
  output        io_Out_enable_valid,
  output        io_Out_enable_bits_control,
  input         io_Out_dataPtrs_field2_0_ready,
  output        io_Out_dataPtrs_field2_0_valid,
  output [63:0] io_Out_dataPtrs_field2_0_bits_data,
  input         io_Out_dataPtrs_field1_0_ready,
  output        io_Out_dataPtrs_field1_0_valid,
  output [63:0] io_Out_dataPtrs_field1_0_bits_data,
  input         io_Out_dataPtrs_field0_0_ready,
  output        io_Out_dataPtrs_field0_0_valid,
  output [63:0] io_Out_dataPtrs_field0_0_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  inputReg_enable_control; // @[SplitDecoupled.scala 220:26]
  reg [63:0] inputReg_dataPtrs_field2_data; // @[SplitDecoupled.scala 220:26]
  reg [63:0] inputReg_dataPtrs_field1_data; // @[SplitDecoupled.scala 220:26]
  reg [63:0] inputReg_dataPtrs_field0_data; // @[SplitDecoupled.scala 220:26]
  reg  enableValidReg; // @[SplitDecoupled.scala 222:31]
  reg  outputPtrsValidReg_0_0; // @[SplitDecoupled.scala 225:53]
  reg  outputPtrsValidReg_1_0; // @[SplitDecoupled.scala 225:53]
  reg  outputPtrsValidReg_2_0; // @[SplitDecoupled.scala 225:53]
  reg  state; // @[SplitDecoupled.scala 260:22]
  wire  _T_1 = ~state; // @[SplitDecoupled.scala 262:24]
  wire  _T_3 = io_In_ready & io_In_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T_3 | state; // @[SplitDecoupled.scala 266:27]
  wire  _GEN_2 = _T_3 | inputReg_enable_control; // @[SplitDecoupled.scala 266:27]
  wire  _T_5 = outputPtrsValidReg_0_0 & outputPtrsValidReg_1_0; // @[SplitDecoupled.scala 247:31]
  wire  _T_6 = _T_5 & outputPtrsValidReg_2_0; // @[SplitDecoupled.scala 247:31]
  wire  _T_7 = ~_T_6; // @[SplitDecoupled.scala 247:7]
  wire  _T_9 = ~enableValidReg; // @[SplitDecoupled.scala 272:43]
  wire  _T_10 = _T_7 & _T_9; // @[SplitDecoupled.scala 272:40]
  wire  _T_12 = io_In_valid & _T_1; // @[SplitDecoupled.scala 280:24]
  wire  _GEN_28 = _T_12 | outputPtrsValidReg_0_0; // @[SplitDecoupled.scala 280:45]
  wire  _T_14 = state & io_Out_dataPtrs_field0_0_ready; // @[SplitDecoupled.scala 283:32]
  wire  _GEN_30 = _T_12 | outputPtrsValidReg_1_0; // @[SplitDecoupled.scala 280:45]
  wire  _T_18 = state & io_Out_dataPtrs_field1_0_ready; // @[SplitDecoupled.scala 283:32]
  wire  _GEN_32 = _T_12 | outputPtrsValidReg_2_0; // @[SplitDecoupled.scala 280:45]
  wire  _T_22 = state & io_Out_dataPtrs_field2_0_ready; // @[SplitDecoupled.scala 283:32]
  wire  _GEN_34 = _T_12 | enableValidReg; // @[SplitDecoupled.scala 305:41]
  wire  _T_26 = state & io_Out_enable_ready; // @[SplitDecoupled.scala 308:28]
  assign io_In_ready = ~state; // @[SplitDecoupled.scala 262:15]
  assign io_Out_enable_valid = enableValidReg; // @[SplitDecoupled.scala 312:23]
  assign io_Out_enable_bits_control = inputReg_enable_control; // @[SplitDecoupled.scala 313:22]
  assign io_Out_dataPtrs_field2_0_valid = outputPtrsValidReg_2_0; // @[SplitDecoupled.scala 286:44]
  assign io_Out_dataPtrs_field2_0_bits_data = inputReg_dataPtrs_field2_data; // @[SplitDecoupled.scala 287:43]
  assign io_Out_dataPtrs_field1_0_valid = outputPtrsValidReg_1_0; // @[SplitDecoupled.scala 286:44]
  assign io_Out_dataPtrs_field1_0_bits_data = inputReg_dataPtrs_field1_data; // @[SplitDecoupled.scala 287:43]
  assign io_Out_dataPtrs_field0_0_valid = outputPtrsValidReg_0_0; // @[SplitDecoupled.scala 286:44]
  assign io_Out_dataPtrs_field0_0_bits_data = inputReg_dataPtrs_field0_data; // @[SplitDecoupled.scala 287:43]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inputReg_enable_control = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  inputReg_dataPtrs_field2_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  inputReg_dataPtrs_field1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  inputReg_dataPtrs_field0_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  enableValidReg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  outputPtrsValidReg_0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  outputPtrsValidReg_1_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  outputPtrsValidReg_2_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      inputReg_enable_control <= 1'h0;
    end else if (_T_1) begin
      inputReg_enable_control <= _GEN_2;
    end
    if (reset) begin
      inputReg_dataPtrs_field2_data <= 64'h0;
    end else if (_T_1) begin
      if (_T_3) begin
        inputReg_dataPtrs_field2_data <= io_In_bits_dataPtrs_field2_data;
      end
    end
    if (reset) begin
      inputReg_dataPtrs_field1_data <= 64'h0;
    end else if (_T_1) begin
      if (_T_3) begin
        inputReg_dataPtrs_field1_data <= io_In_bits_dataPtrs_field1_data;
      end
    end
    if (reset) begin
      inputReg_dataPtrs_field0_data <= 64'h0;
    end else if (_T_1) begin
      if (_T_3) begin
        inputReg_dataPtrs_field0_data <= io_In_bits_dataPtrs_field0_data;
      end
    end
    if (reset) begin
      enableValidReg <= 1'h0;
    end else if (_T_26) begin
      enableValidReg <= 1'h0;
    end else begin
      enableValidReg <= _GEN_34;
    end
    if (reset) begin
      outputPtrsValidReg_0_0 <= 1'h0;
    end else if (_T_14) begin
      outputPtrsValidReg_0_0 <= 1'h0;
    end else begin
      outputPtrsValidReg_0_0 <= _GEN_28;
    end
    if (reset) begin
      outputPtrsValidReg_1_0 <= 1'h0;
    end else if (_T_18) begin
      outputPtrsValidReg_1_0 <= 1'h0;
    end else begin
      outputPtrsValidReg_1_0 <= _GEN_30;
    end
    if (reset) begin
      outputPtrsValidReg_2_0 <= 1'h0;
    end else if (_T_22) begin
      outputPtrsValidReg_2_0 <= 1'h0;
    end else begin
      outputPtrsValidReg_2_0 <= _GEN_32;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_1) begin
      state <= _GEN_0;
    end else if (state) begin
      if (_T_10) begin
        state <= 1'h0;
      end
    end
  end
endmodule
module LoopBlockNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [63:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [63:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [63:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [63:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [63:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [63:0] io_InLiveIn_5_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [63:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field5_1_ready,
  output        io_OutLiveIn_field5_1_valid,
  output [63:0] io_OutLiveIn_field5_1_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [63:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [63:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [63:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [63:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [63:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [63:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [63:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 531:25]
  reg  enable_R_control; // @[LoopBlock.scala 531:25]
  reg  enable_valid_R; // @[LoopBlock.scala 532:31]
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 534:50]
  reg  loop_back_R_0_control; // @[LoopBlock.scala 534:50]
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 535:56]
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 537:54]
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 538:60]
  reg [63:0] in_live_in_R_0_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_1_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_2_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_3_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_4_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_5_data; // @[LoopBlock.scala 540:53]
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 541:59]
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 543:56]
  reg [63:0] in_carry_in_R_0_data; // @[LoopBlock.scala 543:56]
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 544:62]
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_5_1; // @[LoopBlock.scala 556:47]
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_5_1; // @[LoopBlock.scala 560:47]
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 576:44]
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_R_control; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 585:42]
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_R_control; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 588:41]
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 590:47]
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 590:47]
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 591:53]
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 592:52]
  wire  _T_18 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_18 | enable_valid_R; // @[LoopBlock.scala 599:26]
  wire  _T_20 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _GEN_6 = _T_20 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 606:33]
  wire  _GEN_7 = _T_20 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 606:33]
  wire  _GEN_9 = _T_20 | loop_back_valid_R_0; // @[LoopBlock.scala 606:33]
  wire  _T_22 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_22 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 615:35]
  wire  _GEN_13 = _T_22 | loop_finish_valid_R_0; // @[LoopBlock.scala 615:35]
  wire  _T_24 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_24 | in_live_in_valid_R_0; // @[LoopBlock.scala 626:33]
  wire  _T_26 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_26 | in_live_in_valid_R_1; // @[LoopBlock.scala 626:33]
  wire  _T_28 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_25 = _T_28 | in_live_in_valid_R_2; // @[LoopBlock.scala 626:33]
  wire  _T_30 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_30 | in_live_in_valid_R_3; // @[LoopBlock.scala 626:33]
  wire  _T_32 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_33 = _T_32 | in_live_in_valid_R_4; // @[LoopBlock.scala 626:33]
  wire  _T_34 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_37 = _T_34 | in_live_in_valid_R_5; // @[LoopBlock.scala 626:33]
  wire  _T_36 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_41 = _T_36 | in_carry_in_valid_R_0; // @[LoopBlock.scala 644:37]
  wire  _T_37 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_42 = _T_37 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 707:39]
  wire  _T_38 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_43 = _T_38 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 711:38]
  wire  _T_39 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_44 = _T_39 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 716:33]
  wire  _GEN_45 = _T_39 | loop_exit_fire_R_0; // @[LoopBlock.scala 716:33]
  wire  _T_40 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_46 = _T_40 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_47 = _T_40 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _T_41 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_48 = _T_41 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_49 = _T_41 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _T_42 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_50 = _T_42 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_51 = _T_42 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _T_43 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_52 = _T_43 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_53 = _T_43 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _T_44 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_54 = _T_44 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_55 = _T_44 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 725:57]
  wire  _T_45 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_56 = _T_45 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_57 = _T_45 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 725:57]
  wire  _T_46 = io_OutLiveIn_field5_1_ready & io_OutLiveIn_field5_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_58 = _T_46 ? 1'h0 : out_live_in_valid_R_5_1; // @[LoopBlock.scala 725:57]
  wire  _GEN_59 = _T_46 | out_live_in_fire_R_5_1; // @[LoopBlock.scala 725:57]
  wire  _T_47 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_60 = _T_47 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 745:61]
  reg [1:0] state; // @[LoopBlock.scala 864:22]
  wire  _T_51 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_52 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 768:35]
  wire  _T_53 = _T_52 & in_live_in_valid_R_2; // @[LoopBlock.scala 768:35]
  wire  _T_54 = _T_53 & in_live_in_valid_R_3; // @[LoopBlock.scala 768:35]
  wire  _T_55 = _T_54 & in_live_in_valid_R_4; // @[LoopBlock.scala 768:35]
  wire  _T_56 = _T_55 & in_live_in_valid_R_5; // @[LoopBlock.scala 768:35]
  wire  _T_57 = _T_56 & enable_valid_R; // @[LoopBlock.scala 906:28]
  wire  _GEN_62 = enable_R_control | _GEN_46; // @[LoopBlock.scala 907:26]
  wire  _GEN_63 = enable_R_control | _GEN_48; // @[LoopBlock.scala 907:26]
  wire  _GEN_64 = enable_R_control | _GEN_50; // @[LoopBlock.scala 907:26]
  wire  _GEN_65 = enable_R_control | _GEN_52; // @[LoopBlock.scala 907:26]
  wire  _GEN_66 = enable_R_control | _GEN_54; // @[LoopBlock.scala 907:26]
  wire  _GEN_67 = enable_R_control | _GEN_56; // @[LoopBlock.scala 907:26]
  wire  _GEN_68 = enable_R_control | _GEN_58; // @[LoopBlock.scala 907:26]
  wire  _GEN_69 = enable_R_control | _GEN_60; // @[LoopBlock.scala 907:26]
  wire  _GEN_71 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 907:26]
  wire  _GEN_73 = enable_R_control | _GEN_42; // @[LoopBlock.scala 907:26]
  wire  _GEN_77 = enable_R_control | _GEN_43; // @[LoopBlock.scala 907:26]
  wire  _GEN_80 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 907:26]
  wire  _T_61 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_62 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 937:30]
  wire  _T_64 = out_live_in_fire_R_5_0 & out_live_in_fire_R_5_1; // @[LoopBlock.scala 828:65]
  wire  _T_65 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 831:26]
  wire  _T_66 = _T_65 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 831:26]
  wire  _T_67 = _T_66 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 831:26]
  wire  _T_68 = _T_67 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 831:26]
  wire  _T_69 = _T_68 & _T_64; // @[LoopBlock.scala 831:26]
  wire  _T_70 = _T_62 & _T_69; // @[LoopBlock.scala 938:29]
  wire  _T_78 = ~reset; // @[LoopBlock.scala 970:19]
  wire  _GEN_104 = loop_finish_R_0_control | _GEN_44; // @[LoopBlock.scala 974:64]
  wire  _GEN_109 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_112 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_118 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 941:56]
  wire  _GEN_120 = loop_back_R_0_control | _GEN_109; // @[LoopBlock.scala 941:56]
  wire  _GEN_122 = loop_back_R_0_control | _GEN_43; // @[LoopBlock.scala 941:56]
  wire  _GEN_131 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 941:56]
  wire  _GEN_132 = loop_back_R_0_control | _GEN_48; // @[LoopBlock.scala 941:56]
  wire  _GEN_133 = loop_back_R_0_control | _GEN_50; // @[LoopBlock.scala 941:56]
  wire  _GEN_134 = loop_back_R_0_control | _GEN_52; // @[LoopBlock.scala 941:56]
  wire  _GEN_135 = loop_back_R_0_control | _GEN_54; // @[LoopBlock.scala 941:56]
  wire  _GEN_136 = loop_back_R_0_control | _GEN_56; // @[LoopBlock.scala 941:56]
  wire  _GEN_137 = loop_back_R_0_control | _GEN_58; // @[LoopBlock.scala 941:56]
  wire  _GEN_138 = loop_back_R_0_control | _GEN_60; // @[LoopBlock.scala 941:56]
  wire  _T_86 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_399 = ~_T_51; // @[LoopBlock.scala 970:19]
  wire  _GEN_400 = _GEN_399 & _T_61; // @[LoopBlock.scala 970:19]
  wire  _GEN_401 = _GEN_400 & _T_70; // @[LoopBlock.scala 970:19]
  wire  _GEN_402 = _GEN_401 & loop_back_R_0_control; // @[LoopBlock.scala 970:19]
  wire  _GEN_406 = ~loop_back_R_0_control; // @[LoopBlock.scala 988:19]
  wire  _GEN_407 = _GEN_401 & _GEN_406; // @[LoopBlock.scala 988:19]
  wire  _GEN_408 = _GEN_407 & loop_finish_R_0_control; // @[LoopBlock.scala 988:19]
  assign io_enable_ready = ~enable_valid_R; // @[LoopBlock.scala 598:19]
  assign io_InLiveIn_0_ready = ~in_live_in_valid_R_0; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_1_ready = ~in_live_in_valid_R_1; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_2_ready = ~in_live_in_valid_R_2; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_3_ready = ~in_live_in_valid_R_3; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_4_ready = ~in_live_in_valid_R_4; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_5_ready = ~in_live_in_valid_R_5; // @[LoopBlock.scala 625:26]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field5_1_valid = out_live_in_valid_R_5_1; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field5_1_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 667:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 692:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 695:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 694:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 694:30]
  assign io_loopBack_0_ready = ~loop_back_valid_R_0; // @[LoopBlock.scala 605:26]
  assign io_loopFinish_0_ready = ~loop_finish_valid_R_0; // @[LoopBlock.scala 614:28]
  assign io_CarryDepenIn_0_ready = ~in_carry_in_valid_R_0; // @[LoopBlock.scala 643:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 684:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 683:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 683:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 699:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 698:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 698:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  in_live_in_R_3_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  in_live_in_R_4_data = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  in_live_in_R_5_data = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_21[4:0];
  _RAND_22 = {2{`RANDOM}};
  in_carry_in_R_0_data = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  out_live_in_valid_R_5_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  out_live_in_fire_R_5_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  state = _RAND_49[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_51) begin
      if (_T_18) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_61) begin
      if (_T_18) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_18) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_18) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_51) begin
      if (_T_18) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_61) begin
      if (_T_18) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        enable_R_control <= 1'h0;
      end else if (_T_18) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_18) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_51) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_61) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_5;
      end
    end else begin
      enable_valid_R <= _GEN_5;
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else if (_T_51) begin
      if (_T_20) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_taskID <= 5'h0;
        end else if (_T_20) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else if (_T_20) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_taskID <= 5'h0;
      end else if (_T_20) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else begin
      loop_back_R_0_taskID <= _GEN_6;
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else if (_T_51) begin
      if (_T_20) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_control <= 1'h0;
        end else if (_T_20) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else if (_T_20) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_control <= 1'h0;
      end else if (_T_20) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else begin
      loop_back_R_0_control <= _GEN_7;
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else if (_T_51) begin
      loop_back_valid_R_0 <= _GEN_9;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          loop_back_valid_R_0 <= 1'h0;
        end else begin
          loop_back_valid_R_0 <= _GEN_9;
        end
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        loop_back_valid_R_0 <= 1'h0;
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else begin
      loop_back_valid_R_0 <= _GEN_9;
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else if (_T_51) begin
      if (_T_22) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          loop_finish_R_0_control <= 1'h0;
        end else if (_T_22) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else if (_T_22) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_R_0_control <= 1'h0;
      end else if (_T_22) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else begin
      loop_finish_R_0_control <= _GEN_11;
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else if (_T_51) begin
      loop_finish_valid_R_0 <= _GEN_13;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          loop_finish_valid_R_0 <= 1'h0;
        end else begin
          loop_finish_valid_R_0 <= _GEN_13;
        end
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_valid_R_0 <= 1'h0;
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else begin
      loop_finish_valid_R_0 <= _GEN_13;
    end
    if (reset) begin
      in_live_in_R_0_data <= 64'h0;
    end else if (_T_51) begin
      if (_T_24) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_61) begin
      if (_T_24) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_0_data <= 64'h0;
      end else if (_T_24) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_24) begin
      in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
    end
    if (reset) begin
      in_live_in_R_1_data <= 64'h0;
    end else if (_T_51) begin
      if (_T_26) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_61) begin
      if (_T_26) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_1_data <= 64'h0;
      end else if (_T_26) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_26) begin
      in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
    end
    if (reset) begin
      in_live_in_R_2_data <= 64'h0;
    end else if (_T_51) begin
      if (_T_28) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_61) begin
      if (_T_28) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_2_data <= 64'h0;
      end else if (_T_28) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_28) begin
      in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
    end
    if (reset) begin
      in_live_in_R_3_data <= 64'h0;
    end else if (_T_51) begin
      if (_T_30) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_61) begin
      if (_T_30) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_3_data <= 64'h0;
      end else if (_T_30) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_30) begin
      in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
    end
    if (reset) begin
      in_live_in_R_4_data <= 64'h0;
    end else if (_T_51) begin
      if (_T_32) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_61) begin
      if (_T_32) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_4_data <= 64'h0;
      end else if (_T_32) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_32) begin
      in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
    end
    if (reset) begin
      in_live_in_R_5_data <= 64'h0;
    end else if (_T_51) begin
      if (_T_34) begin
        in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
      end
    end else if (_T_61) begin
      if (_T_34) begin
        in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_5_data <= 64'h0;
      end else if (_T_34) begin
        in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
      end
    end else if (_T_34) begin
      in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else if (_T_51) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_61) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_0 <= 1'h0;
      end else begin
        in_live_in_valid_R_0 <= _GEN_17;
      end
    end else begin
      in_live_in_valid_R_0 <= _GEN_17;
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else if (_T_51) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_61) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_1 <= 1'h0;
      end else begin
        in_live_in_valid_R_1 <= _GEN_21;
      end
    end else begin
      in_live_in_valid_R_1 <= _GEN_21;
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else if (_T_51) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_61) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_2 <= 1'h0;
      end else begin
        in_live_in_valid_R_2 <= _GEN_25;
      end
    end else begin
      in_live_in_valid_R_2 <= _GEN_25;
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else if (_T_51) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_61) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_3 <= 1'h0;
      end else begin
        in_live_in_valid_R_3 <= _GEN_29;
      end
    end else begin
      in_live_in_valid_R_3 <= _GEN_29;
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else if (_T_51) begin
      in_live_in_valid_R_4 <= _GEN_33;
    end else if (_T_61) begin
      in_live_in_valid_R_4 <= _GEN_33;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_4 <= 1'h0;
      end else begin
        in_live_in_valid_R_4 <= _GEN_33;
      end
    end else begin
      in_live_in_valid_R_4 <= _GEN_33;
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else if (_T_51) begin
      in_live_in_valid_R_5 <= _GEN_37;
    end else if (_T_61) begin
      in_live_in_valid_R_5 <= _GEN_37;
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_5 <= 1'h0;
      end else begin
        in_live_in_valid_R_5 <= _GEN_37;
      end
    end else begin
      in_live_in_valid_R_5 <= _GEN_37;
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else if (_T_36) begin
      in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
    end
    if (reset) begin
      in_carry_in_R_0_data <= 64'h0;
    end else if (_T_36) begin
      in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else if (_T_51) begin
      in_carry_in_valid_R_0 <= _GEN_41;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          in_carry_in_valid_R_0 <= 1'h0;
        end else begin
          in_carry_in_valid_R_0 <= _GEN_41;
        end
      end else begin
        in_carry_in_valid_R_0 <= _GEN_41;
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        in_carry_in_valid_R_0 <= 1'h0;
      end else begin
        in_carry_in_valid_R_0 <= _GEN_41;
      end
    end else begin
      in_carry_in_valid_R_0 <= _GEN_41;
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_0_0 <= _GEN_62;
      end else if (_T_40) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_0_0 <= _GEN_131;
      end else if (_T_40) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_40) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_1_0 <= _GEN_63;
      end else if (_T_41) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_1_0 <= _GEN_132;
      end else if (_T_41) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_41) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_2_0 <= _GEN_64;
      end else if (_T_42) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_2_0 <= _GEN_133;
      end else if (_T_42) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_42) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_3_0 <= _GEN_65;
      end else if (_T_43) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_3_0 <= _GEN_134;
      end else if (_T_43) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_43) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_4_0 <= _GEN_66;
      end else if (_T_44) begin
        out_live_in_valid_R_4_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_4_0 <= _GEN_135;
      end else if (_T_44) begin
        out_live_in_valid_R_4_0 <= 1'h0;
      end
    end else if (_T_44) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_5_0 <= _GEN_67;
      end else if (_T_45) begin
        out_live_in_valid_R_5_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_5_0 <= _GEN_136;
      end else if (_T_45) begin
        out_live_in_valid_R_5_0 <= 1'h0;
      end
    end else if (_T_45) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_5_1 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_live_in_valid_R_5_1 <= _GEN_68;
      end else if (_T_46) begin
        out_live_in_valid_R_5_1 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_live_in_valid_R_5_1 <= _GEN_137;
      end else if (_T_46) begin
        out_live_in_valid_R_5_1 <= 1'h0;
      end
    end else if (_T_46) begin
      out_live_in_valid_R_5_1 <= 1'h0;
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_0_0 <= _GEN_47;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_0_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_47;
        end
      end else begin
        out_live_in_fire_R_0_0 <= _GEN_47;
      end
    end else begin
      out_live_in_fire_R_0_0 <= _GEN_47;
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_1_0 <= _GEN_49;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_1_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_49;
        end
      end else begin
        out_live_in_fire_R_1_0 <= _GEN_49;
      end
    end else begin
      out_live_in_fire_R_1_0 <= _GEN_49;
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_2_0 <= _GEN_51;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_2_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_51;
        end
      end else begin
        out_live_in_fire_R_2_0 <= _GEN_51;
      end
    end else begin
      out_live_in_fire_R_2_0 <= _GEN_51;
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_3_0 <= _GEN_53;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_3_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_53;
        end
      end else begin
        out_live_in_fire_R_3_0 <= _GEN_53;
      end
    end else begin
      out_live_in_fire_R_3_0 <= _GEN_53;
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_4_0 <= _GEN_55;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_4_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_55;
        end
      end else begin
        out_live_in_fire_R_4_0 <= _GEN_55;
      end
    end else begin
      out_live_in_fire_R_4_0 <= _GEN_55;
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_5_0 <= _GEN_57;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_5_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_57;
        end
      end else begin
        out_live_in_fire_R_5_0 <= _GEN_57;
      end
    end else begin
      out_live_in_fire_R_5_0 <= _GEN_57;
    end
    if (reset) begin
      out_live_in_fire_R_5_1 <= 1'h0;
    end else if (_T_51) begin
      out_live_in_fire_R_5_1 <= _GEN_59;
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_5_1 <= 1'h0;
        end else begin
          out_live_in_fire_R_5_1 <= _GEN_59;
        end
      end else begin
        out_live_in_fire_R_5_1 <= _GEN_59;
      end
    end else begin
      out_live_in_fire_R_5_1 <= _GEN_59;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        out_carry_out_valid_R_0_0 <= _GEN_69;
      end else if (_T_47) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        out_carry_out_valid_R_0_0 <= _GEN_138;
      end else if (_T_47) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_47) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        if (enable_R_control) begin
          active_loop_start_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        active_loop_start_R_control <= _GEN_71;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        active_loop_start_valid_R <= _GEN_73;
      end else if (_T_37) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        active_loop_start_valid_R <= _GEN_118;
      end else if (_T_37) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_37) begin
      active_loop_start_valid_R <= 1'h0;
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        if (enable_R_control) begin
          active_loop_back_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          active_loop_back_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_back_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        if (enable_R_control) begin
          active_loop_back_R_control <= 1'h0;
        end
      end
    end else if (_T_61) begin
      if (_T_70) begin
        active_loop_back_R_control <= _GEN_120;
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        active_loop_back_valid_R <= _GEN_77;
      end else if (_T_38) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        active_loop_back_valid_R <= _GEN_122;
      end else if (_T_38) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_38) begin
      active_loop_back_valid_R <= 1'h0;
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        if (!(enable_R_control)) begin
          loop_exit_R_0_taskID <= 5'h0;
        end
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (!(loop_back_R_0_control)) begin
          if (loop_finish_R_0_control) begin
            loop_exit_R_0_taskID <= loop_back_R_0_taskID;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        loop_exit_R_0_control <= _GEN_80;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (!(loop_back_R_0_control)) begin
          loop_exit_R_0_control <= _GEN_112;
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        if (enable_R_control) begin
          if (_T_39) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= 1'h1;
        end
      end else if (_T_39) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          if (_T_39) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_104;
        end
      end else if (_T_39) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else begin
      loop_exit_valid_R_0 <= _GEN_44;
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_45;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_51) begin
      if (_T_57) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_61) begin
      if (_T_70) begin
        if (loop_back_R_0_control) begin
          state <= 2'h1;
        end else if (loop_finish_R_0_control) begin
          state <= 2'h2;
        end
      end
    end else if (_T_86) begin
      if (loop_exit_fire_R_0) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_402 & _T_78) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_0] [RESTARTED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 970:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_408 & _T_78) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_0] [FIRED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 988:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_408 & _T_78) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_0] [FINAL] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 1003:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [63:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [63:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [63:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [63:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [63:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [63:0] io_InLiveIn_5_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [63:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [63:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field4_1_ready,
  output        io_OutLiveIn_field4_1_valid,
  output [63:0] io_OutLiveIn_field4_1_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [63:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [63:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [63:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [63:0] io_OutLiveIn_field0_0_bits_data,
  input         io_OutLiveIn_field0_1_ready,
  output        io_OutLiveIn_field0_1_valid,
  output [63:0] io_OutLiveIn_field0_1_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [63:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [63:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 531:25]
  reg  enable_R_control; // @[LoopBlock.scala 531:25]
  reg  enable_valid_R; // @[LoopBlock.scala 532:31]
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 534:50]
  reg  loop_back_R_0_control; // @[LoopBlock.scala 534:50]
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 535:56]
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 537:54]
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 538:60]
  reg [63:0] in_live_in_R_0_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_1_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_2_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_3_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_4_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_5_data; // @[LoopBlock.scala 540:53]
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 541:59]
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 543:56]
  reg [63:0] in_carry_in_R_0_data; // @[LoopBlock.scala 543:56]
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 544:62]
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_0_1; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_4_1; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_0_1; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_4_1; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 560:47]
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 576:44]
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_R_control; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 585:42]
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_R_control; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 588:41]
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 590:47]
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 590:47]
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 591:53]
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 592:52]
  wire  _T_18 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_18 | enable_valid_R; // @[LoopBlock.scala 599:26]
  wire  _T_20 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _GEN_6 = _T_20 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 606:33]
  wire  _GEN_7 = _T_20 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 606:33]
  wire  _GEN_9 = _T_20 | loop_back_valid_R_0; // @[LoopBlock.scala 606:33]
  wire  _T_22 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_22 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 615:35]
  wire  _GEN_13 = _T_22 | loop_finish_valid_R_0; // @[LoopBlock.scala 615:35]
  wire  _T_24 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_24 | in_live_in_valid_R_0; // @[LoopBlock.scala 626:33]
  wire  _T_26 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_26 | in_live_in_valid_R_1; // @[LoopBlock.scala 626:33]
  wire  _T_28 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_25 = _T_28 | in_live_in_valid_R_2; // @[LoopBlock.scala 626:33]
  wire  _T_30 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_30 | in_live_in_valid_R_3; // @[LoopBlock.scala 626:33]
  wire  _T_32 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_33 = _T_32 | in_live_in_valid_R_4; // @[LoopBlock.scala 626:33]
  wire  _T_34 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_37 = _T_34 | in_live_in_valid_R_5; // @[LoopBlock.scala 626:33]
  wire  _T_36 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_41 = _T_36 | in_carry_in_valid_R_0; // @[LoopBlock.scala 644:37]
  wire  _T_37 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_42 = _T_37 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 707:39]
  wire  _T_38 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_43 = _T_38 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 711:38]
  wire  _T_39 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_44 = _T_39 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 716:33]
  wire  _GEN_45 = _T_39 | loop_exit_fire_R_0; // @[LoopBlock.scala 716:33]
  wire  _T_40 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_46 = _T_40 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_47 = _T_40 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _T_41 = io_OutLiveIn_field0_1_ready & io_OutLiveIn_field0_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_48 = _T_41 ? 1'h0 : out_live_in_valid_R_0_1; // @[LoopBlock.scala 725:57]
  wire  _GEN_49 = _T_41 | out_live_in_fire_R_0_1; // @[LoopBlock.scala 725:57]
  wire  _T_42 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_50 = _T_42 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_51 = _T_42 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _T_43 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_52 = _T_43 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_53 = _T_43 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _T_44 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_54 = _T_44 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_55 = _T_44 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _T_45 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_56 = _T_45 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_57 = _T_45 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 725:57]
  wire  _T_46 = io_OutLiveIn_field4_1_ready & io_OutLiveIn_field4_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_58 = _T_46 ? 1'h0 : out_live_in_valid_R_4_1; // @[LoopBlock.scala 725:57]
  wire  _GEN_59 = _T_46 | out_live_in_fire_R_4_1; // @[LoopBlock.scala 725:57]
  wire  _T_47 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_60 = _T_47 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_61 = _T_47 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 725:57]
  wire  _T_48 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_62 = _T_48 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 745:61]
  reg [1:0] state; // @[LoopBlock.scala 864:22]
  wire  _T_52 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 768:35]
  wire  _T_54 = _T_53 & in_live_in_valid_R_2; // @[LoopBlock.scala 768:35]
  wire  _T_55 = _T_54 & in_live_in_valid_R_3; // @[LoopBlock.scala 768:35]
  wire  _T_56 = _T_55 & in_live_in_valid_R_4; // @[LoopBlock.scala 768:35]
  wire  _T_57 = _T_56 & in_live_in_valid_R_5; // @[LoopBlock.scala 768:35]
  wire  _T_58 = _T_57 & enable_valid_R; // @[LoopBlock.scala 906:28]
  wire  _GEN_64 = enable_R_control | _GEN_46; // @[LoopBlock.scala 907:26]
  wire  _GEN_65 = enable_R_control | _GEN_48; // @[LoopBlock.scala 907:26]
  wire  _GEN_66 = enable_R_control | _GEN_50; // @[LoopBlock.scala 907:26]
  wire  _GEN_67 = enable_R_control | _GEN_52; // @[LoopBlock.scala 907:26]
  wire  _GEN_68 = enable_R_control | _GEN_54; // @[LoopBlock.scala 907:26]
  wire  _GEN_69 = enable_R_control | _GEN_56; // @[LoopBlock.scala 907:26]
  wire  _GEN_70 = enable_R_control | _GEN_58; // @[LoopBlock.scala 907:26]
  wire  _GEN_71 = enable_R_control | _GEN_60; // @[LoopBlock.scala 907:26]
  wire  _GEN_72 = enable_R_control | _GEN_62; // @[LoopBlock.scala 907:26]
  wire  _GEN_74 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 907:26]
  wire  _GEN_76 = enable_R_control | _GEN_42; // @[LoopBlock.scala 907:26]
  wire  _GEN_80 = enable_R_control | _GEN_43; // @[LoopBlock.scala 907:26]
  wire  _GEN_83 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 907:26]
  wire  _T_62 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_63 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 937:30]
  wire  _T_65 = out_live_in_fire_R_0_0 & out_live_in_fire_R_0_1; // @[LoopBlock.scala 828:65]
  wire  _T_66 = out_live_in_fire_R_4_0 & out_live_in_fire_R_4_1; // @[LoopBlock.scala 828:65]
  wire  _T_67 = _T_65 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 831:26]
  wire  _T_68 = _T_67 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 831:26]
  wire  _T_69 = _T_68 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 831:26]
  wire  _T_70 = _T_69 & _T_66; // @[LoopBlock.scala 831:26]
  wire  _T_71 = _T_70 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 831:26]
  wire  _T_72 = _T_63 & _T_71; // @[LoopBlock.scala 938:29]
  wire  _T_80 = ~reset; // @[LoopBlock.scala 970:19]
  wire  _GEN_108 = loop_finish_R_0_control | _GEN_44; // @[LoopBlock.scala 974:64]
  wire  _GEN_113 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_116 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_122 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 941:56]
  wire  _GEN_124 = loop_back_R_0_control | _GEN_113; // @[LoopBlock.scala 941:56]
  wire  _GEN_126 = loop_back_R_0_control | _GEN_43; // @[LoopBlock.scala 941:56]
  wire  _GEN_136 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 941:56]
  wire  _GEN_137 = loop_back_R_0_control | _GEN_48; // @[LoopBlock.scala 941:56]
  wire  _GEN_138 = loop_back_R_0_control | _GEN_50; // @[LoopBlock.scala 941:56]
  wire  _GEN_139 = loop_back_R_0_control | _GEN_52; // @[LoopBlock.scala 941:56]
  wire  _GEN_140 = loop_back_R_0_control | _GEN_54; // @[LoopBlock.scala 941:56]
  wire  _GEN_141 = loop_back_R_0_control | _GEN_56; // @[LoopBlock.scala 941:56]
  wire  _GEN_142 = loop_back_R_0_control | _GEN_58; // @[LoopBlock.scala 941:56]
  wire  _GEN_143 = loop_back_R_0_control | _GEN_60; // @[LoopBlock.scala 941:56]
  wire  _GEN_144 = loop_back_R_0_control | _GEN_62; // @[LoopBlock.scala 941:56]
  wire  _T_88 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_411 = ~_T_52; // @[LoopBlock.scala 970:19]
  wire  _GEN_412 = _GEN_411 & _T_62; // @[LoopBlock.scala 970:19]
  wire  _GEN_413 = _GEN_412 & _T_72; // @[LoopBlock.scala 970:19]
  wire  _GEN_414 = _GEN_413 & loop_back_R_0_control; // @[LoopBlock.scala 970:19]
  wire  _GEN_418 = ~loop_back_R_0_control; // @[LoopBlock.scala 988:19]
  wire  _GEN_419 = _GEN_413 & _GEN_418; // @[LoopBlock.scala 988:19]
  wire  _GEN_420 = _GEN_419 & loop_finish_R_0_control; // @[LoopBlock.scala 988:19]
  assign io_enable_ready = ~enable_valid_R; // @[LoopBlock.scala 598:19]
  assign io_InLiveIn_0_ready = ~in_live_in_valid_R_0; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_1_ready = ~in_live_in_valid_R_1; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_2_ready = ~in_live_in_valid_R_2; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_3_ready = ~in_live_in_valid_R_3; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_4_ready = ~in_live_in_valid_R_4; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_5_ready = ~in_live_in_valid_R_5; // @[LoopBlock.scala 625:26]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field4_1_valid = out_live_in_valid_R_4_1; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field4_1_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field0_1_valid = out_live_in_valid_R_0_1; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field0_1_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 667:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 692:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 695:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 694:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 694:30]
  assign io_loopBack_0_ready = ~loop_back_valid_R_0; // @[LoopBlock.scala 605:26]
  assign io_loopFinish_0_ready = ~loop_finish_valid_R_0; // @[LoopBlock.scala 614:28]
  assign io_CarryDepenIn_0_ready = ~in_carry_in_valid_R_0; // @[LoopBlock.scala 643:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 684:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 683:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 683:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 699:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 698:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 698:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  in_live_in_R_3_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  in_live_in_R_4_data = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  in_live_in_R_5_data = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_21[4:0];
  _RAND_22 = {2{`RANDOM}};
  in_carry_in_R_0_data = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  out_live_in_valid_R_0_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  out_live_in_valid_R_4_1 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  out_live_in_fire_R_0_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  out_live_in_fire_R_4_1 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  state = _RAND_51[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_52) begin
      if (_T_18) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_62) begin
      if (_T_18) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_18) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_18) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_52) begin
      if (_T_18) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_62) begin
      if (_T_18) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        enable_R_control <= 1'h0;
      end else if (_T_18) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_18) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_52) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_62) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_5;
      end
    end else begin
      enable_valid_R <= _GEN_5;
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else if (_T_52) begin
      if (_T_20) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_taskID <= 5'h0;
        end else if (_T_20) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else if (_T_20) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_taskID <= 5'h0;
      end else if (_T_20) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else begin
      loop_back_R_0_taskID <= _GEN_6;
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else if (_T_52) begin
      if (_T_20) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_control <= 1'h0;
        end else if (_T_20) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else if (_T_20) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_control <= 1'h0;
      end else if (_T_20) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else begin
      loop_back_R_0_control <= _GEN_7;
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else if (_T_52) begin
      loop_back_valid_R_0 <= _GEN_9;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          loop_back_valid_R_0 <= 1'h0;
        end else begin
          loop_back_valid_R_0 <= _GEN_9;
        end
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        loop_back_valid_R_0 <= 1'h0;
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else begin
      loop_back_valid_R_0 <= _GEN_9;
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else if (_T_52) begin
      if (_T_22) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          loop_finish_R_0_control <= 1'h0;
        end else if (_T_22) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else if (_T_22) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_R_0_control <= 1'h0;
      end else if (_T_22) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else begin
      loop_finish_R_0_control <= _GEN_11;
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else if (_T_52) begin
      loop_finish_valid_R_0 <= _GEN_13;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          loop_finish_valid_R_0 <= 1'h0;
        end else begin
          loop_finish_valid_R_0 <= _GEN_13;
        end
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_valid_R_0 <= 1'h0;
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else begin
      loop_finish_valid_R_0 <= _GEN_13;
    end
    if (reset) begin
      in_live_in_R_0_data <= 64'h0;
    end else if (_T_52) begin
      if (_T_24) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_62) begin
      if (_T_24) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_0_data <= 64'h0;
      end else if (_T_24) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_24) begin
      in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
    end
    if (reset) begin
      in_live_in_R_1_data <= 64'h0;
    end else if (_T_52) begin
      if (_T_26) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_62) begin
      if (_T_26) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_1_data <= 64'h0;
      end else if (_T_26) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_26) begin
      in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
    end
    if (reset) begin
      in_live_in_R_2_data <= 64'h0;
    end else if (_T_52) begin
      if (_T_28) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_62) begin
      if (_T_28) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_2_data <= 64'h0;
      end else if (_T_28) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_28) begin
      in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
    end
    if (reset) begin
      in_live_in_R_3_data <= 64'h0;
    end else if (_T_52) begin
      if (_T_30) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_62) begin
      if (_T_30) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_3_data <= 64'h0;
      end else if (_T_30) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_30) begin
      in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
    end
    if (reset) begin
      in_live_in_R_4_data <= 64'h0;
    end else if (_T_52) begin
      if (_T_32) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_62) begin
      if (_T_32) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_4_data <= 64'h0;
      end else if (_T_32) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_32) begin
      in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
    end
    if (reset) begin
      in_live_in_R_5_data <= 64'h0;
    end else if (_T_52) begin
      if (_T_34) begin
        in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
      end
    end else if (_T_62) begin
      if (_T_34) begin
        in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_5_data <= 64'h0;
      end else if (_T_34) begin
        in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
      end
    end else if (_T_34) begin
      in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else if (_T_52) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_62) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_0 <= 1'h0;
      end else begin
        in_live_in_valid_R_0 <= _GEN_17;
      end
    end else begin
      in_live_in_valid_R_0 <= _GEN_17;
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else if (_T_52) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_62) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_1 <= 1'h0;
      end else begin
        in_live_in_valid_R_1 <= _GEN_21;
      end
    end else begin
      in_live_in_valid_R_1 <= _GEN_21;
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else if (_T_52) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_62) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_2 <= 1'h0;
      end else begin
        in_live_in_valid_R_2 <= _GEN_25;
      end
    end else begin
      in_live_in_valid_R_2 <= _GEN_25;
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else if (_T_52) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_62) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_3 <= 1'h0;
      end else begin
        in_live_in_valid_R_3 <= _GEN_29;
      end
    end else begin
      in_live_in_valid_R_3 <= _GEN_29;
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else if (_T_52) begin
      in_live_in_valid_R_4 <= _GEN_33;
    end else if (_T_62) begin
      in_live_in_valid_R_4 <= _GEN_33;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_4 <= 1'h0;
      end else begin
        in_live_in_valid_R_4 <= _GEN_33;
      end
    end else begin
      in_live_in_valid_R_4 <= _GEN_33;
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else if (_T_52) begin
      in_live_in_valid_R_5 <= _GEN_37;
    end else if (_T_62) begin
      in_live_in_valid_R_5 <= _GEN_37;
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_5 <= 1'h0;
      end else begin
        in_live_in_valid_R_5 <= _GEN_37;
      end
    end else begin
      in_live_in_valid_R_5 <= _GEN_37;
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else if (_T_36) begin
      in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
    end
    if (reset) begin
      in_carry_in_R_0_data <= 64'h0;
    end else if (_T_36) begin
      in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else if (_T_52) begin
      in_carry_in_valid_R_0 <= _GEN_41;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          in_carry_in_valid_R_0 <= 1'h0;
        end else begin
          in_carry_in_valid_R_0 <= _GEN_41;
        end
      end else begin
        in_carry_in_valid_R_0 <= _GEN_41;
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        in_carry_in_valid_R_0 <= 1'h0;
      end else begin
        in_carry_in_valid_R_0 <= _GEN_41;
      end
    end else begin
      in_carry_in_valid_R_0 <= _GEN_41;
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_0_0 <= _GEN_64;
      end else if (_T_40) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_0_0 <= _GEN_136;
      end else if (_T_40) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_40) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_0_1 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_0_1 <= _GEN_65;
      end else if (_T_41) begin
        out_live_in_valid_R_0_1 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_0_1 <= _GEN_137;
      end else if (_T_41) begin
        out_live_in_valid_R_0_1 <= 1'h0;
      end
    end else if (_T_41) begin
      out_live_in_valid_R_0_1 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_1_0 <= _GEN_66;
      end else if (_T_42) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_1_0 <= _GEN_138;
      end else if (_T_42) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_42) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_2_0 <= _GEN_67;
      end else if (_T_43) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_2_0 <= _GEN_139;
      end else if (_T_43) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_43) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_3_0 <= _GEN_68;
      end else if (_T_44) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_3_0 <= _GEN_140;
      end else if (_T_44) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_44) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_4_0 <= _GEN_69;
      end else if (_T_45) begin
        out_live_in_valid_R_4_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_4_0 <= _GEN_141;
      end else if (_T_45) begin
        out_live_in_valid_R_4_0 <= 1'h0;
      end
    end else if (_T_45) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_4_1 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_4_1 <= _GEN_70;
      end else if (_T_46) begin
        out_live_in_valid_R_4_1 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_4_1 <= _GEN_142;
      end else if (_T_46) begin
        out_live_in_valid_R_4_1 <= 1'h0;
      end
    end else if (_T_46) begin
      out_live_in_valid_R_4_1 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_live_in_valid_R_5_0 <= _GEN_71;
      end else if (_T_47) begin
        out_live_in_valid_R_5_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_live_in_valid_R_5_0 <= _GEN_143;
      end else if (_T_47) begin
        out_live_in_valid_R_5_0 <= 1'h0;
      end
    end else if (_T_47) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_0_0 <= _GEN_47;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_0_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_47;
        end
      end else begin
        out_live_in_fire_R_0_0 <= _GEN_47;
      end
    end else begin
      out_live_in_fire_R_0_0 <= _GEN_47;
    end
    if (reset) begin
      out_live_in_fire_R_0_1 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_0_1 <= _GEN_49;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_0_1 <= 1'h0;
        end else begin
          out_live_in_fire_R_0_1 <= _GEN_49;
        end
      end else begin
        out_live_in_fire_R_0_1 <= _GEN_49;
      end
    end else begin
      out_live_in_fire_R_0_1 <= _GEN_49;
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_1_0 <= _GEN_51;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_1_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_51;
        end
      end else begin
        out_live_in_fire_R_1_0 <= _GEN_51;
      end
    end else begin
      out_live_in_fire_R_1_0 <= _GEN_51;
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_2_0 <= _GEN_53;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_2_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_53;
        end
      end else begin
        out_live_in_fire_R_2_0 <= _GEN_53;
      end
    end else begin
      out_live_in_fire_R_2_0 <= _GEN_53;
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_3_0 <= _GEN_55;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_3_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_55;
        end
      end else begin
        out_live_in_fire_R_3_0 <= _GEN_55;
      end
    end else begin
      out_live_in_fire_R_3_0 <= _GEN_55;
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_4_0 <= _GEN_57;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_4_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_57;
        end
      end else begin
        out_live_in_fire_R_4_0 <= _GEN_57;
      end
    end else begin
      out_live_in_fire_R_4_0 <= _GEN_57;
    end
    if (reset) begin
      out_live_in_fire_R_4_1 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_4_1 <= _GEN_59;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_4_1 <= 1'h0;
        end else begin
          out_live_in_fire_R_4_1 <= _GEN_59;
        end
      end else begin
        out_live_in_fire_R_4_1 <= _GEN_59;
      end
    end else begin
      out_live_in_fire_R_4_1 <= _GEN_59;
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else if (_T_52) begin
      out_live_in_fire_R_5_0 <= _GEN_61;
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_5_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_61;
        end
      end else begin
        out_live_in_fire_R_5_0 <= _GEN_61;
      end
    end else begin
      out_live_in_fire_R_5_0 <= _GEN_61;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        out_carry_out_valid_R_0_0 <= _GEN_72;
      end else if (_T_48) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        out_carry_out_valid_R_0_0 <= _GEN_144;
      end else if (_T_48) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_48) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        if (enable_R_control) begin
          active_loop_start_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        active_loop_start_R_control <= _GEN_74;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        active_loop_start_valid_R <= _GEN_76;
      end else if (_T_37) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        active_loop_start_valid_R <= _GEN_122;
      end else if (_T_37) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_37) begin
      active_loop_start_valid_R <= 1'h0;
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        if (enable_R_control) begin
          active_loop_back_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          active_loop_back_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_back_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        if (enable_R_control) begin
          active_loop_back_R_control <= 1'h0;
        end
      end
    end else if (_T_62) begin
      if (_T_72) begin
        active_loop_back_R_control <= _GEN_124;
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        active_loop_back_valid_R <= _GEN_80;
      end else if (_T_38) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        active_loop_back_valid_R <= _GEN_126;
      end else if (_T_38) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_38) begin
      active_loop_back_valid_R <= 1'h0;
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        if (!(enable_R_control)) begin
          loop_exit_R_0_taskID <= 5'h0;
        end
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (!(loop_back_R_0_control)) begin
          if (loop_finish_R_0_control) begin
            loop_exit_R_0_taskID <= loop_back_R_0_taskID;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        loop_exit_R_0_control <= _GEN_83;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (!(loop_back_R_0_control)) begin
          loop_exit_R_0_control <= _GEN_116;
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        if (enable_R_control) begin
          if (_T_39) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= 1'h1;
        end
      end else if (_T_39) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          if (_T_39) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_108;
        end
      end else if (_T_39) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else begin
      loop_exit_valid_R_0 <= _GEN_44;
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_45;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_52) begin
      if (_T_58) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_62) begin
      if (_T_72) begin
        if (loop_back_R_0_control) begin
          state <= 2'h1;
        end else if (loop_finish_R_0_control) begin
          state <= 2'h2;
        end
      end
    end else if (_T_88) begin
      if (loop_exit_fire_R_0) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_414 & _T_80) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_1] [RESTARTED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 970:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_420 & _T_80) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_1] [FIRED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 988:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_420 & _T_80) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_1] [FINAL] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 1003:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [63:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [63:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [63:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [63:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [63:0] io_InLiveIn_4_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [63:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [63:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [63:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [63:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [63:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [63:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [63:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 531:25]
  reg  enable_R_control; // @[LoopBlock.scala 531:25]
  reg  enable_valid_R; // @[LoopBlock.scala 532:31]
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 534:50]
  reg  loop_back_R_0_control; // @[LoopBlock.scala 534:50]
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 535:56]
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 537:54]
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 538:60]
  reg [63:0] in_live_in_R_0_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_1_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_2_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_3_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_4_data; // @[LoopBlock.scala 540:53]
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 541:59]
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 543:56]
  reg [63:0] in_carry_in_R_0_data; // @[LoopBlock.scala 543:56]
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 544:62]
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 560:47]
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 576:44]
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_R_control; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 585:42]
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_R_control; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 588:41]
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 590:47]
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 590:47]
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 591:53]
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 592:52]
  wire  _T_17 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_17 | enable_valid_R; // @[LoopBlock.scala 599:26]
  wire  _T_19 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _GEN_6 = _T_19 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 606:33]
  wire  _GEN_7 = _T_19 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 606:33]
  wire  _GEN_9 = _T_19 | loop_back_valid_R_0; // @[LoopBlock.scala 606:33]
  wire  _T_21 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_21 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 615:35]
  wire  _GEN_13 = _T_21 | loop_finish_valid_R_0; // @[LoopBlock.scala 615:35]
  wire  _T_23 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_23 | in_live_in_valid_R_0; // @[LoopBlock.scala 626:33]
  wire  _T_25 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_25 | in_live_in_valid_R_1; // @[LoopBlock.scala 626:33]
  wire  _T_27 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_25 = _T_27 | in_live_in_valid_R_2; // @[LoopBlock.scala 626:33]
  wire  _T_29 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_29 | in_live_in_valid_R_3; // @[LoopBlock.scala 626:33]
  wire  _T_31 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_33 = _T_31 | in_live_in_valid_R_4; // @[LoopBlock.scala 626:33]
  wire  _T_33 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_37 = _T_33 | in_carry_in_valid_R_0; // @[LoopBlock.scala 644:37]
  wire  _T_34 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_38 = _T_34 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 707:39]
  wire  _T_35 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_39 = _T_35 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 711:38]
  wire  _T_36 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_40 = _T_36 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 716:33]
  wire  _GEN_41 = _T_36 | loop_exit_fire_R_0; // @[LoopBlock.scala 716:33]
  wire  _T_37 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_42 = _T_37 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_43 = _T_37 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _T_38 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_44 = _T_38 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_45 = _T_38 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _T_39 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_46 = _T_39 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_47 = _T_39 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _T_40 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_48 = _T_40 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_49 = _T_40 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _T_41 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_50 = _T_41 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_51 = _T_41 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 725:57]
  wire  _T_42 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_52 = _T_42 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 745:61]
  reg [1:0] state; // @[LoopBlock.scala 864:22]
  wire  _T_46 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_47 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 768:35]
  wire  _T_48 = _T_47 & in_live_in_valid_R_2; // @[LoopBlock.scala 768:35]
  wire  _T_49 = _T_48 & in_live_in_valid_R_3; // @[LoopBlock.scala 768:35]
  wire  _T_50 = _T_49 & in_live_in_valid_R_4; // @[LoopBlock.scala 768:35]
  wire  _T_51 = _T_50 & enable_valid_R; // @[LoopBlock.scala 906:28]
  wire  _GEN_54 = enable_R_control | _GEN_42; // @[LoopBlock.scala 907:26]
  wire  _GEN_55 = enable_R_control | _GEN_44; // @[LoopBlock.scala 907:26]
  wire  _GEN_56 = enable_R_control | _GEN_46; // @[LoopBlock.scala 907:26]
  wire  _GEN_57 = enable_R_control | _GEN_48; // @[LoopBlock.scala 907:26]
  wire  _GEN_58 = enable_R_control | _GEN_50; // @[LoopBlock.scala 907:26]
  wire  _GEN_59 = enable_R_control | _GEN_52; // @[LoopBlock.scala 907:26]
  wire  _GEN_61 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 907:26]
  wire  _GEN_63 = enable_R_control | _GEN_38; // @[LoopBlock.scala 907:26]
  wire  _GEN_67 = enable_R_control | _GEN_39; // @[LoopBlock.scala 907:26]
  wire  _GEN_70 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 907:26]
  wire  _T_55 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_56 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 937:30]
  wire  _T_58 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 831:26]
  wire  _T_59 = _T_58 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 831:26]
  wire  _T_60 = _T_59 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 831:26]
  wire  _T_61 = _T_60 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 831:26]
  wire  _T_62 = _T_56 & _T_61; // @[LoopBlock.scala 938:29]
  wire  _T_70 = ~reset; // @[LoopBlock.scala 970:19]
  wire  _GEN_92 = loop_finish_R_0_control | _GEN_40; // @[LoopBlock.scala 974:64]
  wire  _GEN_97 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_100 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_106 = loop_back_R_0_control | _GEN_38; // @[LoopBlock.scala 941:56]
  wire  _GEN_108 = loop_back_R_0_control | _GEN_97; // @[LoopBlock.scala 941:56]
  wire  _GEN_110 = loop_back_R_0_control | _GEN_39; // @[LoopBlock.scala 941:56]
  wire  _GEN_117 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 941:56]
  wire  _GEN_118 = loop_back_R_0_control | _GEN_44; // @[LoopBlock.scala 941:56]
  wire  _GEN_119 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 941:56]
  wire  _GEN_120 = loop_back_R_0_control | _GEN_48; // @[LoopBlock.scala 941:56]
  wire  _GEN_121 = loop_back_R_0_control | _GEN_50; // @[LoopBlock.scala 941:56]
  wire  _GEN_122 = loop_back_R_0_control | _GEN_52; // @[LoopBlock.scala 941:56]
  wire  _T_78 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_355 = ~_T_46; // @[LoopBlock.scala 970:19]
  wire  _GEN_356 = _GEN_355 & _T_55; // @[LoopBlock.scala 970:19]
  wire  _GEN_357 = _GEN_356 & _T_62; // @[LoopBlock.scala 970:19]
  wire  _GEN_358 = _GEN_357 & loop_back_R_0_control; // @[LoopBlock.scala 970:19]
  wire  _GEN_362 = ~loop_back_R_0_control; // @[LoopBlock.scala 988:19]
  wire  _GEN_363 = _GEN_357 & _GEN_362; // @[LoopBlock.scala 988:19]
  wire  _GEN_364 = _GEN_363 & loop_finish_R_0_control; // @[LoopBlock.scala 988:19]
  assign io_enable_ready = ~enable_valid_R; // @[LoopBlock.scala 598:19]
  assign io_InLiveIn_0_ready = ~in_live_in_valid_R_0; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_1_ready = ~in_live_in_valid_R_1; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_2_ready = ~in_live_in_valid_R_2; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_3_ready = ~in_live_in_valid_R_3; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_4_ready = ~in_live_in_valid_R_4; // @[LoopBlock.scala 625:26]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 667:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 692:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 695:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 694:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 694:30]
  assign io_loopBack_0_ready = ~loop_back_valid_R_0; // @[LoopBlock.scala 605:26]
  assign io_loopFinish_0_ready = ~loop_finish_valid_R_0; // @[LoopBlock.scala 614:28]
  assign io_CarryDepenIn_0_ready = ~in_carry_in_valid_R_0; // @[LoopBlock.scala 643:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 684:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 683:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 683:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 699:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 698:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 698:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  in_live_in_R_3_data = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  in_live_in_R_4_data = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_19[4:0];
  _RAND_20 = {2{`RANDOM}};
  in_carry_in_R_0_data = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_33[4:0];
  _RAND_34 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  state = _RAND_43[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_46) begin
      if (_T_17) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_55) begin
      if (_T_17) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_17) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_17) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_46) begin
      if (_T_17) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_55) begin
      if (_T_17) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        enable_R_control <= 1'h0;
      end else if (_T_17) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_17) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_46) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_55) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_5;
      end
    end else begin
      enable_valid_R <= _GEN_5;
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else if (_T_46) begin
      if (_T_19) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_taskID <= 5'h0;
        end else if (_T_19) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else if (_T_19) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_taskID <= 5'h0;
      end else if (_T_19) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else begin
      loop_back_R_0_taskID <= _GEN_6;
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else if (_T_46) begin
      if (_T_19) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_control <= 1'h0;
        end else if (_T_19) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else if (_T_19) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_control <= 1'h0;
      end else if (_T_19) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else begin
      loop_back_R_0_control <= _GEN_7;
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else if (_T_46) begin
      loop_back_valid_R_0 <= _GEN_9;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          loop_back_valid_R_0 <= 1'h0;
        end else begin
          loop_back_valid_R_0 <= _GEN_9;
        end
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        loop_back_valid_R_0 <= 1'h0;
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else begin
      loop_back_valid_R_0 <= _GEN_9;
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else if (_T_46) begin
      if (_T_21) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          loop_finish_R_0_control <= 1'h0;
        end else if (_T_21) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else if (_T_21) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_R_0_control <= 1'h0;
      end else if (_T_21) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else begin
      loop_finish_R_0_control <= _GEN_11;
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else if (_T_46) begin
      loop_finish_valid_R_0 <= _GEN_13;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          loop_finish_valid_R_0 <= 1'h0;
        end else begin
          loop_finish_valid_R_0 <= _GEN_13;
        end
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_valid_R_0 <= 1'h0;
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else begin
      loop_finish_valid_R_0 <= _GEN_13;
    end
    if (reset) begin
      in_live_in_R_0_data <= 64'h0;
    end else if (_T_46) begin
      if (_T_23) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_55) begin
      if (_T_23) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_0_data <= 64'h0;
      end else if (_T_23) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_23) begin
      in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
    end
    if (reset) begin
      in_live_in_R_1_data <= 64'h0;
    end else if (_T_46) begin
      if (_T_25) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_55) begin
      if (_T_25) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_1_data <= 64'h0;
      end else if (_T_25) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_25) begin
      in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
    end
    if (reset) begin
      in_live_in_R_2_data <= 64'h0;
    end else if (_T_46) begin
      if (_T_27) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_55) begin
      if (_T_27) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_2_data <= 64'h0;
      end else if (_T_27) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_27) begin
      in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
    end
    if (reset) begin
      in_live_in_R_3_data <= 64'h0;
    end else if (_T_46) begin
      if (_T_29) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_55) begin
      if (_T_29) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_3_data <= 64'h0;
      end else if (_T_29) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_29) begin
      in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
    end
    if (reset) begin
      in_live_in_R_4_data <= 64'h0;
    end else if (_T_46) begin
      if (_T_31) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_55) begin
      if (_T_31) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_4_data <= 64'h0;
      end else if (_T_31) begin
        in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
      end
    end else if (_T_31) begin
      in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else if (_T_46) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_55) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_0 <= 1'h0;
      end else begin
        in_live_in_valid_R_0 <= _GEN_17;
      end
    end else begin
      in_live_in_valid_R_0 <= _GEN_17;
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else if (_T_46) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_55) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_1 <= 1'h0;
      end else begin
        in_live_in_valid_R_1 <= _GEN_21;
      end
    end else begin
      in_live_in_valid_R_1 <= _GEN_21;
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else if (_T_46) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_55) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_2 <= 1'h0;
      end else begin
        in_live_in_valid_R_2 <= _GEN_25;
      end
    end else begin
      in_live_in_valid_R_2 <= _GEN_25;
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else if (_T_46) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_55) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_3 <= 1'h0;
      end else begin
        in_live_in_valid_R_3 <= _GEN_29;
      end
    end else begin
      in_live_in_valid_R_3 <= _GEN_29;
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else if (_T_46) begin
      in_live_in_valid_R_4 <= _GEN_33;
    end else if (_T_55) begin
      in_live_in_valid_R_4 <= _GEN_33;
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_4 <= 1'h0;
      end else begin
        in_live_in_valid_R_4 <= _GEN_33;
      end
    end else begin
      in_live_in_valid_R_4 <= _GEN_33;
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else if (_T_33) begin
      in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
    end
    if (reset) begin
      in_carry_in_R_0_data <= 64'h0;
    end else if (_T_33) begin
      in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else if (_T_46) begin
      in_carry_in_valid_R_0 <= _GEN_37;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          in_carry_in_valid_R_0 <= 1'h0;
        end else begin
          in_carry_in_valid_R_0 <= _GEN_37;
        end
      end else begin
        in_carry_in_valid_R_0 <= _GEN_37;
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        in_carry_in_valid_R_0 <= 1'h0;
      end else begin
        in_carry_in_valid_R_0 <= _GEN_37;
      end
    end else begin
      in_carry_in_valid_R_0 <= _GEN_37;
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        out_live_in_valid_R_0_0 <= _GEN_54;
      end else if (_T_37) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        out_live_in_valid_R_0_0 <= _GEN_117;
      end else if (_T_37) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_37) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        out_live_in_valid_R_1_0 <= _GEN_55;
      end else if (_T_38) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        out_live_in_valid_R_1_0 <= _GEN_118;
      end else if (_T_38) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_38) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        out_live_in_valid_R_2_0 <= _GEN_56;
      end else if (_T_39) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        out_live_in_valid_R_2_0 <= _GEN_119;
      end else if (_T_39) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_39) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        out_live_in_valid_R_3_0 <= _GEN_57;
      end else if (_T_40) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        out_live_in_valid_R_3_0 <= _GEN_120;
      end else if (_T_40) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_40) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        out_live_in_valid_R_4_0 <= _GEN_58;
      end else if (_T_41) begin
        out_live_in_valid_R_4_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        out_live_in_valid_R_4_0 <= _GEN_121;
      end else if (_T_41) begin
        out_live_in_valid_R_4_0 <= 1'h0;
      end
    end else if (_T_41) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else if (_T_46) begin
      out_live_in_fire_R_0_0 <= _GEN_43;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_0_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_43;
        end
      end else begin
        out_live_in_fire_R_0_0 <= _GEN_43;
      end
    end else begin
      out_live_in_fire_R_0_0 <= _GEN_43;
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else if (_T_46) begin
      out_live_in_fire_R_1_0 <= _GEN_45;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_1_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_45;
        end
      end else begin
        out_live_in_fire_R_1_0 <= _GEN_45;
      end
    end else begin
      out_live_in_fire_R_1_0 <= _GEN_45;
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else if (_T_46) begin
      out_live_in_fire_R_2_0 <= _GEN_47;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_2_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_47;
        end
      end else begin
        out_live_in_fire_R_2_0 <= _GEN_47;
      end
    end else begin
      out_live_in_fire_R_2_0 <= _GEN_47;
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else if (_T_46) begin
      out_live_in_fire_R_3_0 <= _GEN_49;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_3_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_49;
        end
      end else begin
        out_live_in_fire_R_3_0 <= _GEN_49;
      end
    end else begin
      out_live_in_fire_R_3_0 <= _GEN_49;
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else if (_T_46) begin
      out_live_in_fire_R_4_0 <= _GEN_51;
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_4_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_51;
        end
      end else begin
        out_live_in_fire_R_4_0 <= _GEN_51;
      end
    end else begin
      out_live_in_fire_R_4_0 <= _GEN_51;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        out_carry_out_valid_R_0_0 <= _GEN_59;
      end else if (_T_42) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        out_carry_out_valid_R_0_0 <= _GEN_122;
      end else if (_T_42) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_42) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        if (enable_R_control) begin
          active_loop_start_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        active_loop_start_R_control <= _GEN_61;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        active_loop_start_valid_R <= _GEN_63;
      end else if (_T_34) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        active_loop_start_valid_R <= _GEN_106;
      end else if (_T_34) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_34) begin
      active_loop_start_valid_R <= 1'h0;
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        if (enable_R_control) begin
          active_loop_back_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          active_loop_back_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_back_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        if (enable_R_control) begin
          active_loop_back_R_control <= 1'h0;
        end
      end
    end else if (_T_55) begin
      if (_T_62) begin
        active_loop_back_R_control <= _GEN_108;
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        active_loop_back_valid_R <= _GEN_67;
      end else if (_T_35) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        active_loop_back_valid_R <= _GEN_110;
      end else if (_T_35) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_35) begin
      active_loop_back_valid_R <= 1'h0;
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        if (!(enable_R_control)) begin
          loop_exit_R_0_taskID <= 5'h0;
        end
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (!(loop_back_R_0_control)) begin
          if (loop_finish_R_0_control) begin
            loop_exit_R_0_taskID <= loop_back_R_0_taskID;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        loop_exit_R_0_control <= _GEN_70;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (!(loop_back_R_0_control)) begin
          loop_exit_R_0_control <= _GEN_100;
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        if (enable_R_control) begin
          if (_T_36) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= 1'h1;
        end
      end else if (_T_36) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          if (_T_36) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_92;
        end
      end else if (_T_36) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else begin
      loop_exit_valid_R_0 <= _GEN_40;
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_41;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_46) begin
      if (_T_51) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_55) begin
      if (_T_62) begin
        if (loop_back_R_0_control) begin
          state <= 2'h1;
        end else if (loop_finish_R_0_control) begin
          state <= 2'h2;
        end
      end
    end else if (_T_78) begin
      if (loop_exit_fire_R_0) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_358 & _T_70) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_2] [RESTARTED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 970:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_364 & _T_70) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_2] [FIRED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 988:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_364 & _T_70) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_2] [FINAL] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 1003:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [63:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [63:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [63:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [63:0] io_InLiveIn_3_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [63:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [63:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [63:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [63:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [63:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [63:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 531:25]
  reg  enable_R_control; // @[LoopBlock.scala 531:25]
  reg  enable_valid_R; // @[LoopBlock.scala 532:31]
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 534:50]
  reg  loop_back_R_0_control; // @[LoopBlock.scala 534:50]
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 535:56]
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 537:54]
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 538:60]
  reg [63:0] in_live_in_R_0_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_1_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_2_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_3_data; // @[LoopBlock.scala 540:53]
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 541:59]
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 543:56]
  reg [63:0] in_carry_in_R_0_data; // @[LoopBlock.scala 543:56]
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 544:62]
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 560:47]
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 576:44]
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_R_control; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 585:42]
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_R_control; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 588:41]
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 590:47]
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 590:47]
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 591:53]
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 592:52]
  wire  _T_16 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_16 | enable_valid_R; // @[LoopBlock.scala 599:26]
  wire  _T_18 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _GEN_6 = _T_18 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 606:33]
  wire  _GEN_7 = _T_18 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 606:33]
  wire  _GEN_9 = _T_18 | loop_back_valid_R_0; // @[LoopBlock.scala 606:33]
  wire  _T_20 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_20 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 615:35]
  wire  _GEN_13 = _T_20 | loop_finish_valid_R_0; // @[LoopBlock.scala 615:35]
  wire  _T_22 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_22 | in_live_in_valid_R_0; // @[LoopBlock.scala 626:33]
  wire  _T_24 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_24 | in_live_in_valid_R_1; // @[LoopBlock.scala 626:33]
  wire  _T_26 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_25 = _T_26 | in_live_in_valid_R_2; // @[LoopBlock.scala 626:33]
  wire  _T_28 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_28 | in_live_in_valid_R_3; // @[LoopBlock.scala 626:33]
  wire  _T_30 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_33 = _T_30 | in_carry_in_valid_R_0; // @[LoopBlock.scala 644:37]
  wire  _T_31 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_34 = _T_31 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 707:39]
  wire  _T_32 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_35 = _T_32 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 711:38]
  wire  _T_33 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_36 = _T_33 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 716:33]
  wire  _GEN_37 = _T_33 | loop_exit_fire_R_0; // @[LoopBlock.scala 716:33]
  wire  _T_34 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_38 = _T_34 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_39 = _T_34 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _T_35 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_40 = _T_35 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_41 = _T_35 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _T_36 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_42 = _T_36 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_43 = _T_36 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _T_37 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_44 = _T_37 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_45 = _T_37 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 725:57]
  wire  _T_38 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_46 = _T_38 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 745:61]
  reg [1:0] state; // @[LoopBlock.scala 864:22]
  wire  _T_42 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_43 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 768:35]
  wire  _T_44 = _T_43 & in_live_in_valid_R_2; // @[LoopBlock.scala 768:35]
  wire  _T_45 = _T_44 & in_live_in_valid_R_3; // @[LoopBlock.scala 768:35]
  wire  _T_46 = _T_45 & enable_valid_R; // @[LoopBlock.scala 906:28]
  wire  _GEN_48 = enable_R_control | _GEN_38; // @[LoopBlock.scala 907:26]
  wire  _GEN_49 = enable_R_control | _GEN_40; // @[LoopBlock.scala 907:26]
  wire  _GEN_50 = enable_R_control | _GEN_42; // @[LoopBlock.scala 907:26]
  wire  _GEN_51 = enable_R_control | _GEN_44; // @[LoopBlock.scala 907:26]
  wire  _GEN_52 = enable_R_control | _GEN_46; // @[LoopBlock.scala 907:26]
  wire  _GEN_54 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 907:26]
  wire  _GEN_56 = enable_R_control | _GEN_34; // @[LoopBlock.scala 907:26]
  wire  _GEN_60 = enable_R_control | _GEN_35; // @[LoopBlock.scala 907:26]
  wire  _GEN_63 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 907:26]
  wire  _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_51 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 937:30]
  wire  _T_53 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 831:26]
  wire  _T_54 = _T_53 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 831:26]
  wire  _T_55 = _T_54 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 831:26]
  wire  _T_56 = _T_51 & _T_55; // @[LoopBlock.scala 938:29]
  wire  _T_64 = ~reset; // @[LoopBlock.scala 970:19]
  wire  _GEN_84 = loop_finish_R_0_control | _GEN_36; // @[LoopBlock.scala 974:64]
  wire  _GEN_89 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_92 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_98 = loop_back_R_0_control | _GEN_34; // @[LoopBlock.scala 941:56]
  wire  _GEN_100 = loop_back_R_0_control | _GEN_89; // @[LoopBlock.scala 941:56]
  wire  _GEN_102 = loop_back_R_0_control | _GEN_35; // @[LoopBlock.scala 941:56]
  wire  _GEN_108 = loop_back_R_0_control | _GEN_38; // @[LoopBlock.scala 941:56]
  wire  _GEN_109 = loop_back_R_0_control | _GEN_40; // @[LoopBlock.scala 941:56]
  wire  _GEN_110 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 941:56]
  wire  _GEN_111 = loop_back_R_0_control | _GEN_44; // @[LoopBlock.scala 941:56]
  wire  _GEN_112 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 941:56]
  wire  _T_72 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_323 = ~_T_42; // @[LoopBlock.scala 970:19]
  wire  _GEN_324 = _GEN_323 & _T_50; // @[LoopBlock.scala 970:19]
  wire  _GEN_325 = _GEN_324 & _T_56; // @[LoopBlock.scala 970:19]
  wire  _GEN_326 = _GEN_325 & loop_back_R_0_control; // @[LoopBlock.scala 970:19]
  wire  _GEN_330 = ~loop_back_R_0_control; // @[LoopBlock.scala 988:19]
  wire  _GEN_331 = _GEN_325 & _GEN_330; // @[LoopBlock.scala 988:19]
  wire  _GEN_332 = _GEN_331 & loop_finish_R_0_control; // @[LoopBlock.scala 988:19]
  assign io_enable_ready = ~enable_valid_R; // @[LoopBlock.scala 598:19]
  assign io_InLiveIn_0_ready = ~in_live_in_valid_R_0; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_1_ready = ~in_live_in_valid_R_1; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_2_ready = ~in_live_in_valid_R_2; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_3_ready = ~in_live_in_valid_R_3; // @[LoopBlock.scala 625:26]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 667:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 692:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 695:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 694:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 694:30]
  assign io_loopBack_0_ready = ~loop_back_valid_R_0; // @[LoopBlock.scala 605:26]
  assign io_loopFinish_0_ready = ~loop_finish_valid_R_0; // @[LoopBlock.scala 614:28]
  assign io_CarryDepenIn_0_ready = ~in_carry_in_valid_R_0; // @[LoopBlock.scala 643:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 684:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 683:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 683:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 699:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 698:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 698:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  in_live_in_R_3_data = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_17[4:0];
  _RAND_18 = {2{`RANDOM}};
  in_carry_in_R_0_data = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  state = _RAND_39[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_42) begin
      if (_T_16) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_50) begin
      if (_T_16) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_16) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_16) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_42) begin
      if (_T_16) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_50) begin
      if (_T_16) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        enable_R_control <= 1'h0;
      end else if (_T_16) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_16) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_42) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_50) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_5;
      end
    end else begin
      enable_valid_R <= _GEN_5;
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else if (_T_42) begin
      if (_T_18) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_taskID <= 5'h0;
        end else if (_T_18) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else if (_T_18) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_taskID <= 5'h0;
      end else if (_T_18) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else begin
      loop_back_R_0_taskID <= _GEN_6;
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else if (_T_42) begin
      if (_T_18) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_control <= 1'h0;
        end else if (_T_18) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else if (_T_18) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_control <= 1'h0;
      end else if (_T_18) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else begin
      loop_back_R_0_control <= _GEN_7;
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else if (_T_42) begin
      loop_back_valid_R_0 <= _GEN_9;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          loop_back_valid_R_0 <= 1'h0;
        end else begin
          loop_back_valid_R_0 <= _GEN_9;
        end
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        loop_back_valid_R_0 <= 1'h0;
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else begin
      loop_back_valid_R_0 <= _GEN_9;
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else if (_T_42) begin
      if (_T_20) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          loop_finish_R_0_control <= 1'h0;
        end else if (_T_20) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else if (_T_20) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_R_0_control <= 1'h0;
      end else if (_T_20) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else begin
      loop_finish_R_0_control <= _GEN_11;
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else if (_T_42) begin
      loop_finish_valid_R_0 <= _GEN_13;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          loop_finish_valid_R_0 <= 1'h0;
        end else begin
          loop_finish_valid_R_0 <= _GEN_13;
        end
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_valid_R_0 <= 1'h0;
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else begin
      loop_finish_valid_R_0 <= _GEN_13;
    end
    if (reset) begin
      in_live_in_R_0_data <= 64'h0;
    end else if (_T_42) begin
      if (_T_22) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_50) begin
      if (_T_22) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_0_data <= 64'h0;
      end else if (_T_22) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_22) begin
      in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
    end
    if (reset) begin
      in_live_in_R_1_data <= 64'h0;
    end else if (_T_42) begin
      if (_T_24) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_50) begin
      if (_T_24) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_1_data <= 64'h0;
      end else if (_T_24) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_24) begin
      in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
    end
    if (reset) begin
      in_live_in_R_2_data <= 64'h0;
    end else if (_T_42) begin
      if (_T_26) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_50) begin
      if (_T_26) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_2_data <= 64'h0;
      end else if (_T_26) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_26) begin
      in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
    end
    if (reset) begin
      in_live_in_R_3_data <= 64'h0;
    end else if (_T_42) begin
      if (_T_28) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_50) begin
      if (_T_28) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_3_data <= 64'h0;
      end else if (_T_28) begin
        in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
      end
    end else if (_T_28) begin
      in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else if (_T_42) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_50) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_0 <= 1'h0;
      end else begin
        in_live_in_valid_R_0 <= _GEN_17;
      end
    end else begin
      in_live_in_valid_R_0 <= _GEN_17;
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else if (_T_42) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_50) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_1 <= 1'h0;
      end else begin
        in_live_in_valid_R_1 <= _GEN_21;
      end
    end else begin
      in_live_in_valid_R_1 <= _GEN_21;
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else if (_T_42) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_50) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_2 <= 1'h0;
      end else begin
        in_live_in_valid_R_2 <= _GEN_25;
      end
    end else begin
      in_live_in_valid_R_2 <= _GEN_25;
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else if (_T_42) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_50) begin
      in_live_in_valid_R_3 <= _GEN_29;
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_3 <= 1'h0;
      end else begin
        in_live_in_valid_R_3 <= _GEN_29;
      end
    end else begin
      in_live_in_valid_R_3 <= _GEN_29;
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else if (_T_30) begin
      in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
    end
    if (reset) begin
      in_carry_in_R_0_data <= 64'h0;
    end else if (_T_30) begin
      in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else if (_T_42) begin
      in_carry_in_valid_R_0 <= _GEN_33;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          in_carry_in_valid_R_0 <= 1'h0;
        end else begin
          in_carry_in_valid_R_0 <= _GEN_33;
        end
      end else begin
        in_carry_in_valid_R_0 <= _GEN_33;
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        in_carry_in_valid_R_0 <= 1'h0;
      end else begin
        in_carry_in_valid_R_0 <= _GEN_33;
      end
    end else begin
      in_carry_in_valid_R_0 <= _GEN_33;
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        out_live_in_valid_R_0_0 <= _GEN_48;
      end else if (_T_34) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        out_live_in_valid_R_0_0 <= _GEN_108;
      end else if (_T_34) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_34) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        out_live_in_valid_R_1_0 <= _GEN_49;
      end else if (_T_35) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        out_live_in_valid_R_1_0 <= _GEN_109;
      end else if (_T_35) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_35) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        out_live_in_valid_R_2_0 <= _GEN_50;
      end else if (_T_36) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        out_live_in_valid_R_2_0 <= _GEN_110;
      end else if (_T_36) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_36) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        out_live_in_valid_R_3_0 <= _GEN_51;
      end else if (_T_37) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        out_live_in_valid_R_3_0 <= _GEN_111;
      end else if (_T_37) begin
        out_live_in_valid_R_3_0 <= 1'h0;
      end
    end else if (_T_37) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else if (_T_42) begin
      out_live_in_fire_R_0_0 <= _GEN_39;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_0_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_39;
        end
      end else begin
        out_live_in_fire_R_0_0 <= _GEN_39;
      end
    end else begin
      out_live_in_fire_R_0_0 <= _GEN_39;
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else if (_T_42) begin
      out_live_in_fire_R_1_0 <= _GEN_41;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_1_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_41;
        end
      end else begin
        out_live_in_fire_R_1_0 <= _GEN_41;
      end
    end else begin
      out_live_in_fire_R_1_0 <= _GEN_41;
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else if (_T_42) begin
      out_live_in_fire_R_2_0 <= _GEN_43;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_2_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_43;
        end
      end else begin
        out_live_in_fire_R_2_0 <= _GEN_43;
      end
    end else begin
      out_live_in_fire_R_2_0 <= _GEN_43;
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else if (_T_42) begin
      out_live_in_fire_R_3_0 <= _GEN_45;
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_3_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_45;
        end
      end else begin
        out_live_in_fire_R_3_0 <= _GEN_45;
      end
    end else begin
      out_live_in_fire_R_3_0 <= _GEN_45;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        out_carry_out_valid_R_0_0 <= _GEN_52;
      end else if (_T_38) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        out_carry_out_valid_R_0_0 <= _GEN_112;
      end else if (_T_38) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_38) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        if (enable_R_control) begin
          active_loop_start_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        active_loop_start_R_control <= _GEN_54;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        active_loop_start_valid_R <= _GEN_56;
      end else if (_T_31) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        active_loop_start_valid_R <= _GEN_98;
      end else if (_T_31) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_31) begin
      active_loop_start_valid_R <= 1'h0;
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        if (enable_R_control) begin
          active_loop_back_R_taskID <= enable_R_taskID;
        end
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          active_loop_back_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_back_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        if (enable_R_control) begin
          active_loop_back_R_control <= 1'h0;
        end
      end
    end else if (_T_50) begin
      if (_T_56) begin
        active_loop_back_R_control <= _GEN_100;
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        active_loop_back_valid_R <= _GEN_60;
      end else if (_T_32) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        active_loop_back_valid_R <= _GEN_102;
      end else if (_T_32) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_32) begin
      active_loop_back_valid_R <= 1'h0;
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        if (!(enable_R_control)) begin
          loop_exit_R_0_taskID <= 5'h0;
        end
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (!(loop_back_R_0_control)) begin
          if (loop_finish_R_0_control) begin
            loop_exit_R_0_taskID <= loop_back_R_0_taskID;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        loop_exit_R_0_control <= _GEN_63;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (!(loop_back_R_0_control)) begin
          loop_exit_R_0_control <= _GEN_92;
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        if (enable_R_control) begin
          if (_T_33) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= 1'h1;
        end
      end else if (_T_33) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          if (_T_33) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_84;
        end
      end else if (_T_33) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else begin
      loop_exit_valid_R_0 <= _GEN_36;
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_37;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_42) begin
      if (_T_46) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_50) begin
      if (_T_56) begin
        if (loop_back_R_0_control) begin
          state <= 2'h1;
        end else if (loop_finish_R_0_control) begin
          state <= 2'h2;
        end
      end
    end else if (_T_72) begin
      if (loop_exit_fire_R_0) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_326 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_3] [RESTARTED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 970:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_332 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_3] [FIRED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 988:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_332 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_3] [FINAL] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 1003:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [63:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [63:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [63:0] io_InLiveIn_2_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [63:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [63:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [63:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [63:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [63:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  enable_R_control; // @[LoopBlock.scala 531:25]
  reg  enable_valid_R; // @[LoopBlock.scala 532:31]
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 534:50]
  reg  loop_back_R_0_control; // @[LoopBlock.scala 534:50]
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 535:56]
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 537:54]
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 538:60]
  reg [63:0] in_live_in_R_0_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_1_data; // @[LoopBlock.scala 540:53]
  reg [63:0] in_live_in_R_2_data; // @[LoopBlock.scala 540:53]
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 541:59]
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 541:59]
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 543:56]
  reg [63:0] in_carry_in_R_0_data; // @[LoopBlock.scala 543:56]
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 544:62]
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 556:47]
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 560:47]
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 560:47]
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 576:44]
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_R_control; // @[LoopBlock.scala 584:36]
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 585:42]
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_R_control; // @[LoopBlock.scala 587:35]
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 588:41]
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 590:47]
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 590:47]
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 591:53]
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 592:52]
  wire  _T_15 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_15 | enable_valid_R; // @[LoopBlock.scala 599:26]
  wire  _T_17 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  wire [4:0] _GEN_6 = _T_17 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 606:33]
  wire  _GEN_7 = _T_17 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 606:33]
  wire  _GEN_9 = _T_17 | loop_back_valid_R_0; // @[LoopBlock.scala 606:33]
  wire  _T_19 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_19 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 615:35]
  wire  _GEN_13 = _T_19 | loop_finish_valid_R_0; // @[LoopBlock.scala 615:35]
  wire  _T_21 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_21 | in_live_in_valid_R_0; // @[LoopBlock.scala 626:33]
  wire  _T_23 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_23 | in_live_in_valid_R_1; // @[LoopBlock.scala 626:33]
  wire  _T_25 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_25 = _T_25 | in_live_in_valid_R_2; // @[LoopBlock.scala 626:33]
  wire  _T_27 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_27 | in_carry_in_valid_R_0; // @[LoopBlock.scala 644:37]
  wire  _T_28 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_30 = _T_28 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 707:39]
  wire  _T_29 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_31 = _T_29 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 711:38]
  wire  _T_30 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_32 = _T_30 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 716:33]
  wire  _GEN_33 = _T_30 | loop_exit_fire_R_0; // @[LoopBlock.scala 716:33]
  wire  _T_31 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_34 = _T_31 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_35 = _T_31 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 725:57]
  wire  _T_32 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_36 = _T_32 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_37 = _T_32 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 725:57]
  wire  _T_33 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_38 = _T_33 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _GEN_39 = _T_33 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 725:57]
  wire  _T_34 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_40 = _T_34 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 745:61]
  reg [1:0] state; // @[LoopBlock.scala 864:22]
  wire  _T_38 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_39 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 768:35]
  wire  _T_40 = _T_39 & in_live_in_valid_R_2; // @[LoopBlock.scala 768:35]
  wire  _T_41 = _T_40 & enable_valid_R; // @[LoopBlock.scala 906:28]
  wire  _GEN_42 = enable_R_control | _GEN_34; // @[LoopBlock.scala 907:26]
  wire  _GEN_43 = enable_R_control | _GEN_36; // @[LoopBlock.scala 907:26]
  wire  _GEN_44 = enable_R_control | _GEN_38; // @[LoopBlock.scala 907:26]
  wire  _GEN_45 = enable_R_control | _GEN_40; // @[LoopBlock.scala 907:26]
  wire  _GEN_47 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 907:26]
  wire  _GEN_49 = enable_R_control | _GEN_30; // @[LoopBlock.scala 907:26]
  wire  _GEN_53 = enable_R_control | _GEN_31; // @[LoopBlock.scala 907:26]
  wire  _GEN_56 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 907:26]
  wire  _T_45 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_46 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 937:30]
  wire  _T_48 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 831:26]
  wire  _T_49 = _T_48 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 831:26]
  wire  _T_50 = _T_46 & _T_49; // @[LoopBlock.scala 938:29]
  wire  _T_58 = ~reset; // @[LoopBlock.scala 970:19]
  wire  _GEN_76 = loop_finish_R_0_control | _GEN_32; // @[LoopBlock.scala 974:64]
  wire  _GEN_81 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_84 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 974:64]
  wire  _GEN_90 = loop_back_R_0_control | _GEN_30; // @[LoopBlock.scala 941:56]
  wire  _GEN_92 = loop_back_R_0_control | _GEN_81; // @[LoopBlock.scala 941:56]
  wire  _GEN_94 = loop_back_R_0_control | _GEN_31; // @[LoopBlock.scala 941:56]
  wire  _GEN_99 = loop_back_R_0_control | _GEN_34; // @[LoopBlock.scala 941:56]
  wire  _GEN_100 = loop_back_R_0_control | _GEN_36; // @[LoopBlock.scala 941:56]
  wire  _GEN_101 = loop_back_R_0_control | _GEN_38; // @[LoopBlock.scala 941:56]
  wire  _GEN_102 = loop_back_R_0_control | _GEN_40; // @[LoopBlock.scala 941:56]
  wire  _T_66 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _GEN_291 = ~_T_38; // @[LoopBlock.scala 970:19]
  wire  _GEN_292 = _GEN_291 & _T_45; // @[LoopBlock.scala 970:19]
  wire  _GEN_293 = _GEN_292 & _T_50; // @[LoopBlock.scala 970:19]
  wire  _GEN_294 = _GEN_293 & loop_back_R_0_control; // @[LoopBlock.scala 970:19]
  wire  _GEN_298 = ~loop_back_R_0_control; // @[LoopBlock.scala 988:19]
  wire  _GEN_299 = _GEN_293 & _GEN_298; // @[LoopBlock.scala 988:19]
  wire  _GEN_300 = _GEN_299 & loop_finish_R_0_control; // @[LoopBlock.scala 988:19]
  assign io_enable_ready = ~enable_valid_R; // @[LoopBlock.scala 598:19]
  assign io_InLiveIn_0_ready = ~in_live_in_valid_R_0; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_1_ready = ~in_live_in_valid_R_1; // @[LoopBlock.scala 625:26]
  assign io_InLiveIn_2_ready = ~in_live_in_valid_R_2; // @[LoopBlock.scala 625:26]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 667:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 668:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 667:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 692:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 691:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 695:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 694:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 694:30]
  assign io_loopBack_0_ready = ~loop_back_valid_R_0; // @[LoopBlock.scala 605:26]
  assign io_loopFinish_0_ready = ~loop_finish_valid_R_0; // @[LoopBlock.scala 614:28]
  assign io_CarryDepenIn_0_ready = ~in_carry_in_valid_R_0; // @[LoopBlock.scala 643:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 684:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 683:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 683:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 699:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 698:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 698:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  in_live_in_R_0_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  in_live_in_R_1_data = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  in_live_in_R_2_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_14[4:0];
  _RAND_15 = {2{`RANDOM}};
  in_carry_in_R_0_data = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  state = _RAND_34[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_15) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_45) begin
      if (_T_15) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        enable_R_control <= 1'h0;
      end else if (_T_15) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_15) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_38) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_45) begin
      enable_valid_R <= _GEN_5;
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_5;
      end
    end else begin
      enable_valid_R <= _GEN_5;
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_17) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_taskID <= 5'h0;
        end else if (_T_17) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else if (_T_17) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_taskID <= 5'h0;
      end else if (_T_17) begin
        loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
      end
    end else begin
      loop_back_R_0_taskID <= _GEN_6;
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_17) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          loop_back_R_0_control <= 1'h0;
        end else if (_T_17) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else if (_T_17) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        loop_back_R_0_control <= 1'h0;
      end else if (_T_17) begin
        loop_back_R_0_control <= io_loopBack_0_bits_control;
      end
    end else begin
      loop_back_R_0_control <= _GEN_7;
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      loop_back_valid_R_0 <= _GEN_9;
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          loop_back_valid_R_0 <= 1'h0;
        end else begin
          loop_back_valid_R_0 <= _GEN_9;
        end
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        loop_back_valid_R_0 <= 1'h0;
      end else begin
        loop_back_valid_R_0 <= _GEN_9;
      end
    end else begin
      loop_back_valid_R_0 <= _GEN_9;
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_19) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          loop_finish_R_0_control <= 1'h0;
        end else if (_T_19) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else if (_T_19) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_R_0_control <= 1'h0;
      end else if (_T_19) begin
        loop_finish_R_0_control <= io_loopFinish_0_bits_control;
      end
    end else begin
      loop_finish_R_0_control <= _GEN_11;
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      loop_finish_valid_R_0 <= _GEN_13;
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          loop_finish_valid_R_0 <= 1'h0;
        end else begin
          loop_finish_valid_R_0 <= _GEN_13;
        end
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        loop_finish_valid_R_0 <= 1'h0;
      end else begin
        loop_finish_valid_R_0 <= _GEN_13;
      end
    end else begin
      loop_finish_valid_R_0 <= _GEN_13;
    end
    if (reset) begin
      in_live_in_R_0_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_21) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_45) begin
      if (_T_21) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_0_data <= 64'h0;
      end else if (_T_21) begin
        in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
      end
    end else if (_T_21) begin
      in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
    end
    if (reset) begin
      in_live_in_R_1_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_23) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_45) begin
      if (_T_23) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_1_data <= 64'h0;
      end else if (_T_23) begin
        in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
      end
    end else if (_T_23) begin
      in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
    end
    if (reset) begin
      in_live_in_R_2_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_25) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_45) begin
      if (_T_25) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_R_2_data <= 64'h0;
      end else if (_T_25) begin
        in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
      end
    end else if (_T_25) begin
      in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_45) begin
      in_live_in_valid_R_0 <= _GEN_17;
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_0 <= 1'h0;
      end else begin
        in_live_in_valid_R_0 <= _GEN_17;
      end
    end else begin
      in_live_in_valid_R_0 <= _GEN_17;
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else if (_T_38) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_45) begin
      in_live_in_valid_R_1 <= _GEN_21;
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_1 <= 1'h0;
      end else begin
        in_live_in_valid_R_1 <= _GEN_21;
      end
    end else begin
      in_live_in_valid_R_1 <= _GEN_21;
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else if (_T_38) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_45) begin
      in_live_in_valid_R_2 <= _GEN_25;
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_live_in_valid_R_2 <= 1'h0;
      end else begin
        in_live_in_valid_R_2 <= _GEN_25;
      end
    end else begin
      in_live_in_valid_R_2 <= _GEN_25;
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else if (_T_27) begin
      in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
    end
    if (reset) begin
      in_carry_in_R_0_data <= 64'h0;
    end else if (_T_27) begin
      in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      in_carry_in_valid_R_0 <= _GEN_29;
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          in_carry_in_valid_R_0 <= 1'h0;
        end else begin
          in_carry_in_valid_R_0 <= _GEN_29;
        end
      end else begin
        in_carry_in_valid_R_0 <= _GEN_29;
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        in_carry_in_valid_R_0 <= 1'h0;
      end else begin
        in_carry_in_valid_R_0 <= _GEN_29;
      end
    end else begin
      in_carry_in_valid_R_0 <= _GEN_29;
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        out_live_in_valid_R_0_0 <= _GEN_42;
      end else if (_T_31) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        out_live_in_valid_R_0_0 <= _GEN_99;
      end else if (_T_31) begin
        out_live_in_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_31) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        out_live_in_valid_R_1_0 <= _GEN_43;
      end else if (_T_32) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        out_live_in_valid_R_1_0 <= _GEN_100;
      end else if (_T_32) begin
        out_live_in_valid_R_1_0 <= 1'h0;
      end
    end else if (_T_32) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        out_live_in_valid_R_2_0 <= _GEN_44;
      end else if (_T_33) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        out_live_in_valid_R_2_0 <= _GEN_101;
      end else if (_T_33) begin
        out_live_in_valid_R_2_0 <= 1'h0;
      end
    end else if (_T_33) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else if (_T_38) begin
      out_live_in_fire_R_0_0 <= _GEN_35;
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_0_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_35;
        end
      end else begin
        out_live_in_fire_R_0_0 <= _GEN_35;
      end
    end else begin
      out_live_in_fire_R_0_0 <= _GEN_35;
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else if (_T_38) begin
      out_live_in_fire_R_1_0 <= _GEN_37;
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_1_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_37;
        end
      end else begin
        out_live_in_fire_R_1_0 <= _GEN_37;
      end
    end else begin
      out_live_in_fire_R_1_0 <= _GEN_37;
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else if (_T_38) begin
      out_live_in_fire_R_2_0 <= _GEN_39;
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          out_live_in_fire_R_2_0 <= 1'h0;
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_39;
        end
      end else begin
        out_live_in_fire_R_2_0 <= _GEN_39;
      end
    end else begin
      out_live_in_fire_R_2_0 <= _GEN_39;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        out_carry_out_valid_R_0_0 <= _GEN_45;
      end else if (_T_34) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        out_carry_out_valid_R_0_0 <= _GEN_102;
      end else if (_T_34) begin
        out_carry_out_valid_R_0_0 <= 1'h0;
      end
    end else if (_T_34) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        if (enable_R_control) begin
          active_loop_start_R_taskID <= 5'h0;
        end
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        active_loop_start_R_control <= _GEN_47;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end else if (loop_finish_R_0_control) begin
          active_loop_start_R_control <= 1'h0;
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        active_loop_start_valid_R <= _GEN_49;
      end else if (_T_28) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        active_loop_start_valid_R <= _GEN_90;
      end else if (_T_28) begin
        active_loop_start_valid_R <= 1'h0;
      end
    end else if (_T_28) begin
      active_loop_start_valid_R <= 1'h0;
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        if (enable_R_control) begin
          active_loop_back_R_taskID <= 5'h0;
        end
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          active_loop_back_R_taskID <= loop_back_R_0_taskID;
        end else if (loop_finish_R_0_control) begin
          active_loop_back_R_taskID <= 5'h0;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        if (enable_R_control) begin
          active_loop_back_R_control <= 1'h0;
        end
      end
    end else if (_T_45) begin
      if (_T_50) begin
        active_loop_back_R_control <= _GEN_92;
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        active_loop_back_valid_R <= _GEN_53;
      end else if (_T_29) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        active_loop_back_valid_R <= _GEN_94;
      end else if (_T_29) begin
        active_loop_back_valid_R <= 1'h0;
      end
    end else if (_T_29) begin
      active_loop_back_valid_R <= 1'h0;
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        if (!(enable_R_control)) begin
          loop_exit_R_0_taskID <= 5'h0;
        end
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (!(loop_back_R_0_control)) begin
          if (loop_finish_R_0_control) begin
            loop_exit_R_0_taskID <= loop_back_R_0_taskID;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        loop_exit_R_0_control <= _GEN_56;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (!(loop_back_R_0_control)) begin
          loop_exit_R_0_control <= _GEN_84;
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        if (enable_R_control) begin
          if (_T_30) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= 1'h1;
        end
      end else if (_T_30) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          if (_T_30) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_76;
        end
      end else if (_T_30) begin
        loop_exit_valid_R_0 <= 1'h0;
      end
    end else begin
      loop_exit_valid_R_0 <= _GEN_32;
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_33;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_38) begin
      if (_T_41) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_45) begin
      if (_T_50) begin
        if (loop_back_R_0_control) begin
          state <= 2'h1;
        end else if (loop_finish_R_0_control) begin
          state <= 2'h2;
        end
      end
    end else if (_T_66) begin
      if (loop_exit_fire_R_0) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_294 & _T_58) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_4] [RESTARTED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 970:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & _T_58) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_4] [FIRED] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 988:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_300 & _T_58) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOOP] [Loop_4] [FINAL] [Cycle: %d]\n",io_activate_loop_start_bits_taskID,cycleCount); // @[LoopBlock.scala 1003:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode(
  input   clock,
  input   reset,
  output  io_predicateIn_0_ready,
  input   io_predicateIn_0_valid,
  input   io_predicateIn_0_bits_control,
  input   io_Out_0_ready,
  output  io_Out_0_valid,
  output  io_Out_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  in_data_R_0_control; // @[BasicBlock.scala 224:46]
  reg  in_data_valid_R_0; // @[BasicBlock.scala 225:52]
  reg  output_valid_R_0; // @[BasicBlock.scala 228:49]
  reg  output_fire_R_0; // @[BasicBlock.scala 229:48]
  wire  _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 234:36]
  wire  _GEN_5 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 234:36]
  wire  _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 246:28]
  wire  out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 258:85]
  reg  state; // @[BasicBlock.scala 289:22]
  wire  _T_15 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_19 = ~reset; // @[BasicBlock.scala 311:17]
  wire  _GEN_8 = _GEN_5 | output_valid_R_0; // @[BasicBlock.scala 301:9]
  wire  _GEN_10 = _GEN_5 | state; // @[BasicBlock.scala 301:9]
  wire  _GEN_31 = _T_15 & _GEN_5; // @[BasicBlock.scala 311:17]
  assign io_predicateIn_0_ready = ~in_data_valid_R_0; // @[BasicBlock.scala 233:29]
  assign io_Out_0_valid = _T_15 ? _GEN_8 : output_valid_R_0; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else if (_T_15) begin
      if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (state) begin
      if (out_fire_mask_0) begin
        in_data_R_0_control <= 1'h0;
      end else if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (_T_7) begin
      in_data_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      in_data_valid_R_0 <= _GEN_5;
    end else if (state) begin
      if (out_fire_mask_0) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_5;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_5;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      if (_GEN_5) begin
        output_valid_R_0 <= _T_17;
      end else if (_T_8) begin
        output_valid_R_0 <= 1'h0;
      end
    end else if (_T_8) begin
      output_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else if (_T_15) begin
      output_fire_R_0 <= _GEN_6;
    end else if (state) begin
      if (out_fire_mask_0) begin
        output_fire_R_0 <= 1'h0;
      end else begin
        output_fire_R_0 <= _GEN_6;
      end
    end else begin
      output_fire_R_0 <= _GEN_6;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_15) begin
      state <= _GEN_10;
    end else if (state) begin
      if (out_fire_mask_0) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] [bb_entry0] [Out: %d] [Cycle: %d]\n",5'h0,_GEN_3,cycleCount); // @[BasicBlock.scala 311:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  out_ready_R_0; // @[HandShaking.scala 780:28]
  reg  out_ready_R_1; // @[HandShaking.scala 780:28]
  reg  out_ready_R_2; // @[HandShaking.scala 780:28]
  reg  out_valid_R_0; // @[HandShaking.scala 781:28]
  reg  out_valid_R_1; // @[HandShaking.scala 781:28]
  reg  out_valid_R_2; // @[HandShaking.scala 781:28]
  reg  mask_valid_R_0; // @[HandShaking.scala 785:46]
  wire  _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 794:29]
  wire  _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 794:29]
  wire  _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 794:29]
  wire  _T_5 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_5 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 805:32]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_9 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 65:51]
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 65:51]
  reg  predicate_control_R_0; // @[BasicBlock.scala 66:36]
  reg  predicate_control_R_1; // @[BasicBlock.scala 66:36]
  reg  predicate_valid_R_0; // @[BasicBlock.scala 67:54]
  reg  predicate_valid_R_1; // @[BasicBlock.scala 67:54]
  reg  state; // @[BasicBlock.scala 70:22]
  wire  predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 76:58]
  wire [4:0] predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 77:62]
  wire  _T_13 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = _T_13 | predicate_valid_R_0; // @[BasicBlock.scala 80:91]
  wire  _T_16 = _T_14 | predicate_valid_R_1; // @[BasicBlock.scala 80:91]
  wire  start = _T_15 & _T_16; // @[BasicBlock.scala 80:107]
  wire [1:0] _T_21 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:52]
  wire  _T_22 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_20 = start | _GEN_1; // @[BasicBlock.scala 115:19]
  wire  _GEN_21 = start | _GEN_3; // @[BasicBlock.scala 115:19]
  wire  _GEN_22 = start | _GEN_5; // @[BasicBlock.scala 115:19]
  wire  _GEN_23 = start | _GEN_7; // @[BasicBlock.scala 115:19]
  wire  _GEN_24 = start | state; // @[BasicBlock.scala 115:19]
  wire [2:0] _T_26 = {out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 834:17]
  wire  _T_27 = &_T_26; // @[HandShaking.scala 834:24]
  wire  _T_31 = ~reset; // @[BasicBlock.scala 129:19]
  wire  _GEN_50 = ~_T_22; // @[BasicBlock.scala 129:19]
  wire  _GEN_51 = _GEN_50 & state; // @[BasicBlock.scala 129:19]
  wire  _GEN_52 = _GEN_51 & _T_27; // @[BasicBlock.scala 129:19]
  wire  _GEN_53 = _GEN_52 & predicate; // @[BasicBlock.scala 129:19]
  wire  _GEN_57 = ~predicate; // @[BasicBlock.scala 134:19]
  wire  _GEN_58 = _GEN_52 & _GEN_57; // @[BasicBlock.scala 134:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 804:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 793:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 793:21]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 793:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_predicateIn_0_ready = ~predicate_valid_R_0; // @[BasicBlock.scala 88:29]
  assign io_predicateIn_1_ready = ~predicate_valid_R_1; // @[BasicBlock.scala 88:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_27) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_2) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_27) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_3) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (state) begin
      if (_T_27) begin
        out_ready_R_2 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (_T_4) begin
      out_ready_R_2 <= io_Out_2_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      out_valid_R_0 <= _GEN_20;
    end else if (_T_2) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_22) begin
      out_valid_R_1 <= _GEN_21;
    end else if (_T_3) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_22) begin
      out_valid_R_2 <= _GEN_22;
    end else if (_T_4) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      mask_valid_R_0 <= _GEN_23;
    end else if (_T_5) begin
      mask_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_9;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else if (_T_13) begin
      predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else if (_T_13) begin
      predicate_in_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else if (_T_14) begin
      predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else if (_T_14) begin
      predicate_in_R_1_control <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else if (_T_13) begin
      predicate_control_R_0 <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else if (_T_14) begin
      predicate_control_R_1 <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      predicate_valid_R_0 <= _T_15;
    end else if (state) begin
      if (_T_27) begin
        predicate_valid_R_0 <= 1'h0;
      end else begin
        predicate_valid_R_0 <= _T_15;
      end
    end else begin
      predicate_valid_R_0 <= _T_15;
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else if (_T_22) begin
      predicate_valid_R_1 <= _T_16;
    end else if (state) begin
      if (_T_27) begin
        predicate_valid_R_1 <= 1'h0;
      end else begin
        predicate_valid_R_1 <= _T_16;
      end
    end else begin
      predicate_valid_R_1 <= _T_16;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_27) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_31) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] bb_loopkk1] [Mask: 0x%x]\n",predicate_task,_T_21); // @[BasicBlock.scala 129:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_58 & _T_31) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] bb_loopkk1: Output fired @ %d -> 0 predicate\n",cycleCount); // @[BasicBlock.scala 134:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_1(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  out_ready_R_0; // @[HandShaking.scala 780:28]
  reg  out_ready_R_1; // @[HandShaking.scala 780:28]
  reg  out_ready_R_2; // @[HandShaking.scala 780:28]
  reg  out_valid_R_0; // @[HandShaking.scala 781:28]
  reg  out_valid_R_1; // @[HandShaking.scala 781:28]
  reg  out_valid_R_2; // @[HandShaking.scala 781:28]
  reg  mask_valid_R_0; // @[HandShaking.scala 785:46]
  wire  _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 794:29]
  wire  _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 794:29]
  wire  _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 794:29]
  wire  _T_5 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_5 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 805:32]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_9 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 65:51]
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 65:51]
  reg  predicate_control_R_0; // @[BasicBlock.scala 66:36]
  reg  predicate_control_R_1; // @[BasicBlock.scala 66:36]
  reg  predicate_valid_R_0; // @[BasicBlock.scala 67:54]
  reg  predicate_valid_R_1; // @[BasicBlock.scala 67:54]
  reg  state; // @[BasicBlock.scala 70:22]
  wire  predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 76:58]
  wire [4:0] predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 77:62]
  wire  _T_13 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_15 = _T_13 | predicate_valid_R_0; // @[BasicBlock.scala 80:91]
  wire  _T_16 = _T_14 | predicate_valid_R_1; // @[BasicBlock.scala 80:91]
  wire  start = _T_15 & _T_16; // @[BasicBlock.scala 80:107]
  wire [1:0] _T_21 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:52]
  wire  _T_22 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_20 = start | _GEN_1; // @[BasicBlock.scala 115:19]
  wire  _GEN_21 = start | _GEN_3; // @[BasicBlock.scala 115:19]
  wire  _GEN_22 = start | _GEN_5; // @[BasicBlock.scala 115:19]
  wire  _GEN_23 = start | _GEN_7; // @[BasicBlock.scala 115:19]
  wire  _GEN_24 = start | state; // @[BasicBlock.scala 115:19]
  wire [2:0] _T_26 = {out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 834:17]
  wire  _T_27 = &_T_26; // @[HandShaking.scala 834:24]
  wire  _T_31 = ~reset; // @[BasicBlock.scala 129:19]
  wire  _GEN_50 = ~_T_22; // @[BasicBlock.scala 129:19]
  wire  _GEN_51 = _GEN_50 & state; // @[BasicBlock.scala 129:19]
  wire  _GEN_52 = _GEN_51 & _T_27; // @[BasicBlock.scala 129:19]
  wire  _GEN_53 = _GEN_52 & predicate; // @[BasicBlock.scala 129:19]
  wire  _GEN_57 = ~predicate; // @[BasicBlock.scala 134:19]
  wire  _GEN_58 = _GEN_52 & _GEN_57; // @[BasicBlock.scala 134:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 804:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 793:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 793:21]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 793:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_predicateIn_0_ready = ~predicate_valid_R_0; // @[BasicBlock.scala 88:29]
  assign io_predicateIn_1_ready = ~predicate_valid_R_1; // @[BasicBlock.scala 88:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_27) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_2) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_27) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_3) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (state) begin
      if (_T_27) begin
        out_ready_R_2 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (_T_4) begin
      out_ready_R_2 <= io_Out_2_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      out_valid_R_0 <= _GEN_20;
    end else if (_T_2) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_22) begin
      out_valid_R_1 <= _GEN_21;
    end else if (_T_3) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_22) begin
      out_valid_R_2 <= _GEN_22;
    end else if (_T_4) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      mask_valid_R_0 <= _GEN_23;
    end else if (_T_5) begin
      mask_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_9;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else if (_T_13) begin
      predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else if (_T_13) begin
      predicate_in_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else if (_T_14) begin
      predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else if (_T_14) begin
      predicate_in_R_1_control <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else if (_T_13) begin
      predicate_control_R_0 <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else if (_T_14) begin
      predicate_control_R_1 <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      predicate_valid_R_0 <= _T_15;
    end else if (state) begin
      if (_T_27) begin
        predicate_valid_R_0 <= 1'h0;
      end else begin
        predicate_valid_R_0 <= _T_15;
      end
    end else begin
      predicate_valid_R_0 <= _T_15;
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else if (_T_22) begin
      predicate_valid_R_1 <= _T_16;
    end else if (state) begin
      if (_T_27) begin
        predicate_valid_R_1 <= 1'h0;
      end else begin
        predicate_valid_R_1 <= _T_16;
      end
    end else begin
      predicate_valid_R_1 <= _T_16;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_27) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_31) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] bb_loopi2] [Mask: 0x%x]\n",predicate_task,_T_21); // @[BasicBlock.scala 129:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_58 & _T_31) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] bb_loopi2: Output fired @ %d -> 0 predicate\n",cycleCount); // @[BasicBlock.scala 134:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_2(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg  out_ready_R_0; // @[HandShaking.scala 780:28]
  reg  out_ready_R_1; // @[HandShaking.scala 780:28]
  reg  out_ready_R_2; // @[HandShaking.scala 780:28]
  reg  out_ready_R_3; // @[HandShaking.scala 780:28]
  reg  out_ready_R_4; // @[HandShaking.scala 780:28]
  reg  out_valid_R_0; // @[HandShaking.scala 781:28]
  reg  out_valid_R_1; // @[HandShaking.scala 781:28]
  reg  out_valid_R_2; // @[HandShaking.scala 781:28]
  reg  out_valid_R_3; // @[HandShaking.scala 781:28]
  reg  out_valid_R_4; // @[HandShaking.scala 781:28]
  reg  mask_valid_R_0; // @[HandShaking.scala 785:46]
  wire  _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 794:29]
  wire  _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 794:29]
  wire  _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 794:29]
  wire  _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 794:29]
  wire  _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 794:29]
  wire  _T_7 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_7 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 805:32]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_11 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 65:51]
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 65:51]
  reg  predicate_control_R_0; // @[BasicBlock.scala 66:36]
  reg  predicate_control_R_1; // @[BasicBlock.scala 66:36]
  reg  predicate_valid_R_0; // @[BasicBlock.scala 67:54]
  reg  predicate_valid_R_1; // @[BasicBlock.scala 67:54]
  reg  state; // @[BasicBlock.scala 70:22]
  wire  predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 76:58]
  wire [4:0] predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 77:62]
  wire  _T_15 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_16 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_17 = _T_15 | predicate_valid_R_0; // @[BasicBlock.scala 80:91]
  wire  _T_18 = _T_16 | predicate_valid_R_1; // @[BasicBlock.scala 80:91]
  wire  start = _T_17 & _T_18; // @[BasicBlock.scala 80:107]
  wire [1:0] _T_23 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:52]
  wire  _T_24 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_24 = start | _GEN_1; // @[BasicBlock.scala 115:19]
  wire  _GEN_25 = start | _GEN_3; // @[BasicBlock.scala 115:19]
  wire  _GEN_26 = start | _GEN_5; // @[BasicBlock.scala 115:19]
  wire  _GEN_27 = start | _GEN_7; // @[BasicBlock.scala 115:19]
  wire  _GEN_28 = start | _GEN_9; // @[BasicBlock.scala 115:19]
  wire  _GEN_29 = start | _GEN_11; // @[BasicBlock.scala 115:19]
  wire  _GEN_30 = start | state; // @[BasicBlock.scala 115:19]
  wire [4:0] _T_30 = {out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 834:17]
  wire  _T_31 = &_T_30; // @[HandShaking.scala 834:24]
  wire  _T_35 = ~reset; // @[BasicBlock.scala 129:19]
  wire  _GEN_64 = ~_T_24; // @[BasicBlock.scala 129:19]
  wire  _GEN_65 = _GEN_64 & state; // @[BasicBlock.scala 129:19]
  wire  _GEN_66 = _GEN_65 & _T_31; // @[BasicBlock.scala 129:19]
  wire  _GEN_67 = _GEN_66 & predicate; // @[BasicBlock.scala 129:19]
  wire  _GEN_71 = ~predicate; // @[BasicBlock.scala 134:19]
  wire  _GEN_72 = _GEN_66 & _GEN_71; // @[BasicBlock.scala 134:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 804:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 793:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 793:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 793:21]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 793:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 793:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_predicateIn_0_ready = ~predicate_valid_R_0; // @[BasicBlock.scala 88:29]
  assign io_predicateIn_1_ready = ~predicate_valid_R_1; // @[BasicBlock.scala 88:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cycleCount = _RAND_11[14:0];
  _RAND_12 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  state = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_24) begin
      if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_31) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_2) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_24) begin
      if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_31) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_3) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else if (_T_24) begin
      if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (state) begin
      if (_T_31) begin
        out_ready_R_2 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (_T_4) begin
      out_ready_R_2 <= io_Out_2_ready;
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else if (_T_24) begin
      if (_T_5) begin
        out_ready_R_3 <= io_Out_3_ready;
      end
    end else if (state) begin
      if (_T_31) begin
        out_ready_R_3 <= 1'h0;
      end else if (_T_5) begin
        out_ready_R_3 <= io_Out_3_ready;
      end
    end else if (_T_5) begin
      out_ready_R_3 <= io_Out_3_ready;
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else if (_T_24) begin
      if (_T_6) begin
        out_ready_R_4 <= io_Out_4_ready;
      end
    end else if (state) begin
      if (_T_31) begin
        out_ready_R_4 <= 1'h0;
      end else if (_T_6) begin
        out_ready_R_4 <= io_Out_4_ready;
      end
    end else if (_T_6) begin
      out_ready_R_4 <= io_Out_4_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_24) begin
      out_valid_R_0 <= _GEN_24;
    end else if (_T_2) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_24) begin
      out_valid_R_1 <= _GEN_25;
    end else if (_T_3) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_24) begin
      out_valid_R_2 <= _GEN_26;
    end else if (_T_4) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else if (_T_24) begin
      out_valid_R_3 <= _GEN_27;
    end else if (_T_5) begin
      out_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else if (_T_24) begin
      out_valid_R_4 <= _GEN_28;
    end else if (_T_6) begin
      out_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else if (_T_24) begin
      mask_valid_R_0 <= _GEN_29;
    end else if (_T_7) begin
      mask_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_11;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else if (_T_15) begin
      predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else if (_T_15) begin
      predicate_in_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else if (_T_16) begin
      predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else if (_T_16) begin
      predicate_in_R_1_control <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else if (_T_15) begin
      predicate_control_R_0 <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else if (_T_16) begin
      predicate_control_R_1 <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else if (_T_24) begin
      predicate_valid_R_0 <= _T_17;
    end else if (state) begin
      if (_T_31) begin
        predicate_valid_R_0 <= 1'h0;
      end else begin
        predicate_valid_R_0 <= _T_17;
      end
    end else begin
      predicate_valid_R_0 <= _T_17;
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else if (_T_24) begin
      predicate_valid_R_1 <= _T_18;
    end else if (state) begin
      if (_T_31) begin
        predicate_valid_R_1 <= 1'h0;
      end else begin
        predicate_valid_R_1 <= _T_18;
      end
    end else begin
      predicate_valid_R_1 <= _T_18;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_24) begin
      state <= _GEN_30;
    end else if (state) begin
      if (_T_31) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_35) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] bb_loopk3] [Mask: 0x%x]\n",predicate_task,_T_23); // @[BasicBlock.scala 129:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_72 & _T_35) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] bb_loopk3: Output fired @ %d -> 0 predicate\n",cycleCount); // @[BasicBlock.scala 134:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_3(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg  out_ready_R_0; // @[HandShaking.scala 780:28]
  reg  out_ready_R_1; // @[HandShaking.scala 780:28]
  reg  out_ready_R_2; // @[HandShaking.scala 780:28]
  reg  out_ready_R_3; // @[HandShaking.scala 780:28]
  reg  out_ready_R_4; // @[HandShaking.scala 780:28]
  reg  out_ready_R_5; // @[HandShaking.scala 780:28]
  reg  out_ready_R_6; // @[HandShaking.scala 780:28]
  reg  out_ready_R_7; // @[HandShaking.scala 780:28]
  reg  out_ready_R_8; // @[HandShaking.scala 780:28]
  reg  out_ready_R_9; // @[HandShaking.scala 780:28]
  reg  out_valid_R_0; // @[HandShaking.scala 781:28]
  reg  out_valid_R_1; // @[HandShaking.scala 781:28]
  reg  out_valid_R_2; // @[HandShaking.scala 781:28]
  reg  out_valid_R_3; // @[HandShaking.scala 781:28]
  reg  out_valid_R_4; // @[HandShaking.scala 781:28]
  reg  out_valid_R_5; // @[HandShaking.scala 781:28]
  reg  out_valid_R_6; // @[HandShaking.scala 781:28]
  reg  out_valid_R_7; // @[HandShaking.scala 781:28]
  reg  out_valid_R_8; // @[HandShaking.scala 781:28]
  reg  out_valid_R_9; // @[HandShaking.scala 781:28]
  reg  mask_valid_R_0; // @[HandShaking.scala 785:46]
  wire  _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 794:29]
  wire  _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 794:29]
  wire  _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 794:29]
  wire  _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 794:29]
  wire  _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 794:29]
  wire  _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 794:29]
  wire  _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 794:29]
  wire  _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 794:29]
  wire  _T_10 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_10 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 794:29]
  wire  _T_11 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_19 = _T_11 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 794:29]
  wire  _T_12 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_12 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 805:32]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_16 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 65:51]
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 65:51]
  reg  predicate_control_R_0; // @[BasicBlock.scala 66:36]
  reg  predicate_control_R_1; // @[BasicBlock.scala 66:36]
  reg  predicate_valid_R_0; // @[BasicBlock.scala 67:54]
  reg  predicate_valid_R_1; // @[BasicBlock.scala 67:54]
  reg  state; // @[BasicBlock.scala 70:22]
  wire  predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 76:58]
  wire [4:0] predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 77:62]
  wire  _T_20 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_21 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_22 = _T_20 | predicate_valid_R_0; // @[BasicBlock.scala 80:91]
  wire  _T_23 = _T_21 | predicate_valid_R_1; // @[BasicBlock.scala 80:91]
  wire  start = _T_22 & _T_23; // @[BasicBlock.scala 80:107]
  wire [1:0] _T_28 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:52]
  wire  _T_29 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_34 = start | _GEN_1; // @[BasicBlock.scala 115:19]
  wire  _GEN_35 = start | _GEN_3; // @[BasicBlock.scala 115:19]
  wire  _GEN_36 = start | _GEN_5; // @[BasicBlock.scala 115:19]
  wire  _GEN_37 = start | _GEN_7; // @[BasicBlock.scala 115:19]
  wire  _GEN_38 = start | _GEN_9; // @[BasicBlock.scala 115:19]
  wire  _GEN_39 = start | _GEN_11; // @[BasicBlock.scala 115:19]
  wire  _GEN_40 = start | _GEN_13; // @[BasicBlock.scala 115:19]
  wire  _GEN_41 = start | _GEN_15; // @[BasicBlock.scala 115:19]
  wire  _GEN_42 = start | _GEN_17; // @[BasicBlock.scala 115:19]
  wire  _GEN_43 = start | _GEN_19; // @[BasicBlock.scala 115:19]
  wire  _GEN_44 = start | _GEN_21; // @[BasicBlock.scala 115:19]
  wire  _GEN_45 = start | state; // @[BasicBlock.scala 115:19]
  wire [9:0] _T_40 = {out_ready_R_9,out_ready_R_8,out_ready_R_7,out_ready_R_6,out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 834:17]
  wire  _T_41 = &_T_40; // @[HandShaking.scala 834:24]
  wire  _T_45 = ~reset; // @[BasicBlock.scala 129:19]
  wire  _GEN_99 = ~_T_29; // @[BasicBlock.scala 129:19]
  wire  _GEN_100 = _GEN_99 & state; // @[BasicBlock.scala 129:19]
  wire  _GEN_101 = _GEN_100 & _T_41; // @[BasicBlock.scala 129:19]
  wire  _GEN_102 = _GEN_101 & predicate; // @[BasicBlock.scala 129:19]
  wire  _GEN_106 = ~predicate; // @[BasicBlock.scala 134:19]
  wire  _GEN_107 = _GEN_101 & _GEN_106; // @[BasicBlock.scala 134:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 804:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 793:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 793:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 793:21]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 793:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 793:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 793:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 793:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 793:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 793:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_8_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 793:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_9_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_predicateIn_0_ready = ~predicate_valid_R_0; // @[BasicBlock.scala 88:29]
  assign io_predicateIn_1_ready = ~predicate_valid_R_1; // @[BasicBlock.scala 88:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  cycleCount = _RAND_21[14:0];
  _RAND_22 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  state = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_29) begin
      if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_2) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_29) begin
      if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_3) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else if (_T_29) begin
      if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_2 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (_T_4) begin
      out_ready_R_2 <= io_Out_2_ready;
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else if (_T_29) begin
      if (_T_5) begin
        out_ready_R_3 <= io_Out_3_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_3 <= 1'h0;
      end else if (_T_5) begin
        out_ready_R_3 <= io_Out_3_ready;
      end
    end else if (_T_5) begin
      out_ready_R_3 <= io_Out_3_ready;
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else if (_T_29) begin
      if (_T_6) begin
        out_ready_R_4 <= io_Out_4_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_4 <= 1'h0;
      end else if (_T_6) begin
        out_ready_R_4 <= io_Out_4_ready;
      end
    end else if (_T_6) begin
      out_ready_R_4 <= io_Out_4_ready;
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else if (_T_29) begin
      if (_T_7) begin
        out_ready_R_5 <= io_Out_5_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_5 <= 1'h0;
      end else if (_T_7) begin
        out_ready_R_5 <= io_Out_5_ready;
      end
    end else if (_T_7) begin
      out_ready_R_5 <= io_Out_5_ready;
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else if (_T_29) begin
      if (_T_8) begin
        out_ready_R_6 <= io_Out_6_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_6 <= 1'h0;
      end else if (_T_8) begin
        out_ready_R_6 <= io_Out_6_ready;
      end
    end else if (_T_8) begin
      out_ready_R_6 <= io_Out_6_ready;
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else if (_T_29) begin
      if (_T_9) begin
        out_ready_R_7 <= io_Out_7_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_7 <= 1'h0;
      end else if (_T_9) begin
        out_ready_R_7 <= io_Out_7_ready;
      end
    end else if (_T_9) begin
      out_ready_R_7 <= io_Out_7_ready;
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else if (_T_29) begin
      if (_T_10) begin
        out_ready_R_8 <= io_Out_8_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_8 <= 1'h0;
      end else if (_T_10) begin
        out_ready_R_8 <= io_Out_8_ready;
      end
    end else if (_T_10) begin
      out_ready_R_8 <= io_Out_8_ready;
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else if (_T_29) begin
      if (_T_11) begin
        out_ready_R_9 <= io_Out_9_ready;
      end
    end else if (state) begin
      if (_T_41) begin
        out_ready_R_9 <= 1'h0;
      end else if (_T_11) begin
        out_ready_R_9 <= io_Out_9_ready;
      end
    end else if (_T_11) begin
      out_ready_R_9 <= io_Out_9_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_0 <= _GEN_34;
    end else if (_T_2) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_1 <= _GEN_35;
    end else if (_T_3) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_2 <= _GEN_36;
    end else if (_T_4) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_3 <= _GEN_37;
    end else if (_T_5) begin
      out_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_4 <= _GEN_38;
    end else if (_T_6) begin
      out_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_5 <= _GEN_39;
    end else if (_T_7) begin
      out_valid_R_5 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_6 <= _GEN_40;
    end else if (_T_8) begin
      out_valid_R_6 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_7 <= _GEN_41;
    end else if (_T_9) begin
      out_valid_R_7 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_8 <= _GEN_42;
    end else if (_T_10) begin
      out_valid_R_8 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else if (_T_29) begin
      out_valid_R_9 <= _GEN_43;
    end else if (_T_11) begin
      out_valid_R_9 <= 1'h0;
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else if (_T_29) begin
      mask_valid_R_0 <= _GEN_44;
    end else if (_T_12) begin
      mask_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_16;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else if (_T_20) begin
      predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else if (_T_20) begin
      predicate_in_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else if (_T_21) begin
      predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else if (_T_21) begin
      predicate_in_R_1_control <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else if (_T_20) begin
      predicate_control_R_0 <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else if (_T_21) begin
      predicate_control_R_1 <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else if (_T_29) begin
      predicate_valid_R_0 <= _T_22;
    end else if (state) begin
      if (_T_41) begin
        predicate_valid_R_0 <= 1'h0;
      end else begin
        predicate_valid_R_0 <= _T_22;
      end
    end else begin
      predicate_valid_R_0 <= _T_22;
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else if (_T_29) begin
      predicate_valid_R_1 <= _T_23;
    end else if (state) begin
      if (_T_41) begin
        predicate_valid_R_1 <= 1'h0;
      end else begin
        predicate_valid_R_1 <= _T_23;
      end
    end else begin
      predicate_valid_R_1 <= _T_23;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_29) begin
      state <= _GEN_45;
    end else if (state) begin
      if (_T_41) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_102 & _T_45) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] bb_for_body94] [Mask: 0x%x]\n",predicate_task,_T_28); // @[BasicBlock.scala 129:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_107 & _T_45) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] bb_for_body94: Output fired @ %d -> 0 predicate\n",cycleCount); // @[BasicBlock.scala 134:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_4(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output [4:0] io_Out_10_bits_taskID,
  output       io_Out_10_bits_control,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output [4:0] io_Out_11_bits_taskID,
  output       io_Out_11_bits_control,
  input        io_Out_12_ready,
  output       io_Out_12_valid,
  output [4:0] io_Out_12_bits_taskID,
  output       io_Out_12_bits_control,
  input        io_Out_13_ready,
  output       io_Out_13_valid,
  output [4:0] io_Out_13_bits_taskID,
  output       io_Out_13_bits_control,
  input        io_Out_14_ready,
  output       io_Out_14_valid,
  output [4:0] io_Out_14_bits_taskID,
  output       io_Out_14_bits_control,
  input        io_Out_15_ready,
  output       io_Out_15_valid,
  output [4:0] io_Out_15_bits_taskID,
  output       io_Out_15_bits_control,
  input        io_Out_16_ready,
  output       io_Out_16_valid,
  output [4:0] io_Out_16_bits_taskID,
  output       io_Out_16_bits_control,
  input        io_Out_17_ready,
  output       io_Out_17_valid,
  output [4:0] io_Out_17_bits_taskID,
  output       io_Out_17_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
`endif // RANDOMIZE_REG_INIT
  reg  out_ready_R_0; // @[HandShaking.scala 780:28]
  reg  out_ready_R_1; // @[HandShaking.scala 780:28]
  reg  out_ready_R_2; // @[HandShaking.scala 780:28]
  reg  out_ready_R_3; // @[HandShaking.scala 780:28]
  reg  out_ready_R_4; // @[HandShaking.scala 780:28]
  reg  out_ready_R_5; // @[HandShaking.scala 780:28]
  reg  out_ready_R_6; // @[HandShaking.scala 780:28]
  reg  out_ready_R_7; // @[HandShaking.scala 780:28]
  reg  out_ready_R_8; // @[HandShaking.scala 780:28]
  reg  out_ready_R_9; // @[HandShaking.scala 780:28]
  reg  out_ready_R_10; // @[HandShaking.scala 780:28]
  reg  out_ready_R_11; // @[HandShaking.scala 780:28]
  reg  out_ready_R_12; // @[HandShaking.scala 780:28]
  reg  out_ready_R_13; // @[HandShaking.scala 780:28]
  reg  out_ready_R_14; // @[HandShaking.scala 780:28]
  reg  out_ready_R_15; // @[HandShaking.scala 780:28]
  reg  out_ready_R_16; // @[HandShaking.scala 780:28]
  reg  out_ready_R_17; // @[HandShaking.scala 780:28]
  reg  out_valid_R_0; // @[HandShaking.scala 781:28]
  reg  out_valid_R_1; // @[HandShaking.scala 781:28]
  reg  out_valid_R_2; // @[HandShaking.scala 781:28]
  reg  out_valid_R_3; // @[HandShaking.scala 781:28]
  reg  out_valid_R_4; // @[HandShaking.scala 781:28]
  reg  out_valid_R_5; // @[HandShaking.scala 781:28]
  reg  out_valid_R_6; // @[HandShaking.scala 781:28]
  reg  out_valid_R_7; // @[HandShaking.scala 781:28]
  reg  out_valid_R_8; // @[HandShaking.scala 781:28]
  reg  out_valid_R_9; // @[HandShaking.scala 781:28]
  reg  out_valid_R_10; // @[HandShaking.scala 781:28]
  reg  out_valid_R_11; // @[HandShaking.scala 781:28]
  reg  out_valid_R_12; // @[HandShaking.scala 781:28]
  reg  out_valid_R_13; // @[HandShaking.scala 781:28]
  reg  out_valid_R_14; // @[HandShaking.scala 781:28]
  reg  out_valid_R_15; // @[HandShaking.scala 781:28]
  reg  out_valid_R_16; // @[HandShaking.scala 781:28]
  reg  out_valid_R_17; // @[HandShaking.scala 781:28]
  reg  mask_valid_R_0; // @[HandShaking.scala 785:46]
  wire  _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 794:29]
  wire  _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 794:29]
  wire  _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 794:29]
  wire  _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 794:29]
  wire  _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 794:29]
  wire  _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 794:29]
  wire  _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 794:29]
  wire  _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 794:29]
  wire  _T_10 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_10 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 794:29]
  wire  _T_11 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_19 = _T_11 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 794:29]
  wire  _T_12 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_21 = _T_12 ? 1'h0 : out_valid_R_10; // @[HandShaking.scala 794:29]
  wire  _T_13 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_23 = _T_13 ? 1'h0 : out_valid_R_11; // @[HandShaking.scala 794:29]
  wire  _T_14 = io_Out_12_ready & io_Out_12_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_25 = _T_14 ? 1'h0 : out_valid_R_12; // @[HandShaking.scala 794:29]
  wire  _T_15 = io_Out_13_ready & io_Out_13_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_27 = _T_15 ? 1'h0 : out_valid_R_13; // @[HandShaking.scala 794:29]
  wire  _T_16 = io_Out_14_ready & io_Out_14_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_29 = _T_16 ? 1'h0 : out_valid_R_14; // @[HandShaking.scala 794:29]
  wire  _T_17 = io_Out_15_ready & io_Out_15_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_31 = _T_17 ? 1'h0 : out_valid_R_15; // @[HandShaking.scala 794:29]
  wire  _T_18 = io_Out_16_ready & io_Out_16_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_33 = _T_18 ? 1'h0 : out_valid_R_16; // @[HandShaking.scala 794:29]
  wire  _T_19 = io_Out_17_ready & io_Out_17_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_35 = _T_19 ? 1'h0 : out_valid_R_17; // @[HandShaking.scala 794:29]
  wire  _T_20 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_37 = _T_20 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 805:32]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_24 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 65:51]
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 65:51]
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 65:51]
  reg  predicate_control_R_0; // @[BasicBlock.scala 66:36]
  reg  predicate_control_R_1; // @[BasicBlock.scala 66:36]
  reg  predicate_valid_R_0; // @[BasicBlock.scala 67:54]
  reg  predicate_valid_R_1; // @[BasicBlock.scala 67:54]
  reg  state; // @[BasicBlock.scala 70:22]
  wire  predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 76:58]
  wire [4:0] predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 77:62]
  wire  _T_28 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_29 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = _T_28 | predicate_valid_R_0; // @[BasicBlock.scala 80:91]
  wire  _T_31 = _T_29 | predicate_valid_R_1; // @[BasicBlock.scala 80:91]
  wire  start = _T_30 & _T_31; // @[BasicBlock.scala 80:107]
  wire [1:0] _T_36 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:52]
  wire  _T_37 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_50 = start | _GEN_1; // @[BasicBlock.scala 115:19]
  wire  _GEN_51 = start | _GEN_3; // @[BasicBlock.scala 115:19]
  wire  _GEN_52 = start | _GEN_5; // @[BasicBlock.scala 115:19]
  wire  _GEN_53 = start | _GEN_7; // @[BasicBlock.scala 115:19]
  wire  _GEN_54 = start | _GEN_9; // @[BasicBlock.scala 115:19]
  wire  _GEN_55 = start | _GEN_11; // @[BasicBlock.scala 115:19]
  wire  _GEN_56 = start | _GEN_13; // @[BasicBlock.scala 115:19]
  wire  _GEN_57 = start | _GEN_15; // @[BasicBlock.scala 115:19]
  wire  _GEN_58 = start | _GEN_17; // @[BasicBlock.scala 115:19]
  wire  _GEN_59 = start | _GEN_19; // @[BasicBlock.scala 115:19]
  wire  _GEN_60 = start | _GEN_21; // @[BasicBlock.scala 115:19]
  wire  _GEN_61 = start | _GEN_23; // @[BasicBlock.scala 115:19]
  wire  _GEN_62 = start | _GEN_25; // @[BasicBlock.scala 115:19]
  wire  _GEN_63 = start | _GEN_27; // @[BasicBlock.scala 115:19]
  wire  _GEN_64 = start | _GEN_29; // @[BasicBlock.scala 115:19]
  wire  _GEN_65 = start | _GEN_31; // @[BasicBlock.scala 115:19]
  wire  _GEN_66 = start | _GEN_33; // @[BasicBlock.scala 115:19]
  wire  _GEN_67 = start | _GEN_35; // @[BasicBlock.scala 115:19]
  wire  _GEN_68 = start | _GEN_37; // @[BasicBlock.scala 115:19]
  wire  _GEN_69 = start | state; // @[BasicBlock.scala 115:19]
  wire [8:0] _T_47 = {out_ready_R_8,out_ready_R_7,out_ready_R_6,out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 834:17]
  wire [17:0] _T_56 = {out_ready_R_17,out_ready_R_16,out_ready_R_15,out_ready_R_14,out_ready_R_13,out_ready_R_12,out_ready_R_11,out_ready_R_10,out_ready_R_9,_T_47}; // @[HandShaking.scala 834:17]
  wire  _T_57 = &_T_56; // @[HandShaking.scala 834:24]
  wire  _T_61 = ~reset; // @[BasicBlock.scala 129:19]
  wire  _GEN_155 = ~_T_37; // @[BasicBlock.scala 129:19]
  wire  _GEN_156 = _GEN_155 & state; // @[BasicBlock.scala 129:19]
  wire  _GEN_157 = _GEN_156 & _T_57; // @[BasicBlock.scala 129:19]
  wire  _GEN_158 = _GEN_157 & predicate; // @[BasicBlock.scala 129:19]
  wire  _GEN_162 = ~predicate; // @[BasicBlock.scala 134:19]
  wire  _GEN_163 = _GEN_157 & _GEN_162; // @[BasicBlock.scala 134:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 804:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 105:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 793:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 793:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 793:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 793:21]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 793:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 793:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 793:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 793:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 793:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_8_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 793:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_9_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_10_valid = out_valid_R_10; // @[HandShaking.scala 793:21]
  assign io_Out_10_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_10_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_11_valid = out_valid_R_11; // @[HandShaking.scala 793:21]
  assign io_Out_11_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_11_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_12_valid = out_valid_R_12; // @[HandShaking.scala 793:21]
  assign io_Out_12_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_12_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_13_valid = out_valid_R_13; // @[HandShaking.scala 793:21]
  assign io_Out_13_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_13_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_14_valid = out_valid_R_14; // @[HandShaking.scala 793:21]
  assign io_Out_14_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_14_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_15_valid = out_valid_R_15; // @[HandShaking.scala 793:21]
  assign io_Out_15_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_15_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_16_valid = out_valid_R_16; // @[HandShaking.scala 793:21]
  assign io_Out_16_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_16_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_Out_17_valid = out_valid_R_17; // @[HandShaking.scala 793:21]
  assign io_Out_17_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 99:27]
  assign io_Out_17_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 98:28]
  assign io_predicateIn_0_ready = ~predicate_valid_R_0; // @[BasicBlock.scala 88:29]
  assign io_predicateIn_1_ready = ~predicate_valid_R_1; // @[BasicBlock.scala 88:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_ready_R_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  out_ready_R_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  out_ready_R_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  out_ready_R_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  out_ready_R_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  out_ready_R_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  out_valid_R_10 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  out_valid_R_11 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  out_valid_R_12 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  out_valid_R_13 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  out_valid_R_14 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  out_valid_R_15 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  out_valid_R_16 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  out_valid_R_17 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  cycleCount = _RAND_37[14:0];
  _RAND_38 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  state = _RAND_46[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_37) begin
      if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_2) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_37) begin
      if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_3) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_3) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else if (_T_37) begin
      if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_2 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_2 <= io_Out_2_ready;
      end
    end else if (_T_4) begin
      out_ready_R_2 <= io_Out_2_ready;
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else if (_T_37) begin
      if (_T_5) begin
        out_ready_R_3 <= io_Out_3_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_3 <= 1'h0;
      end else if (_T_5) begin
        out_ready_R_3 <= io_Out_3_ready;
      end
    end else if (_T_5) begin
      out_ready_R_3 <= io_Out_3_ready;
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else if (_T_37) begin
      if (_T_6) begin
        out_ready_R_4 <= io_Out_4_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_4 <= 1'h0;
      end else if (_T_6) begin
        out_ready_R_4 <= io_Out_4_ready;
      end
    end else if (_T_6) begin
      out_ready_R_4 <= io_Out_4_ready;
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else if (_T_37) begin
      if (_T_7) begin
        out_ready_R_5 <= io_Out_5_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_5 <= 1'h0;
      end else if (_T_7) begin
        out_ready_R_5 <= io_Out_5_ready;
      end
    end else if (_T_7) begin
      out_ready_R_5 <= io_Out_5_ready;
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else if (_T_37) begin
      if (_T_8) begin
        out_ready_R_6 <= io_Out_6_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_6 <= 1'h0;
      end else if (_T_8) begin
        out_ready_R_6 <= io_Out_6_ready;
      end
    end else if (_T_8) begin
      out_ready_R_6 <= io_Out_6_ready;
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else if (_T_37) begin
      if (_T_9) begin
        out_ready_R_7 <= io_Out_7_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_7 <= 1'h0;
      end else if (_T_9) begin
        out_ready_R_7 <= io_Out_7_ready;
      end
    end else if (_T_9) begin
      out_ready_R_7 <= io_Out_7_ready;
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else if (_T_37) begin
      if (_T_10) begin
        out_ready_R_8 <= io_Out_8_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_8 <= 1'h0;
      end else if (_T_10) begin
        out_ready_R_8 <= io_Out_8_ready;
      end
    end else if (_T_10) begin
      out_ready_R_8 <= io_Out_8_ready;
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else if (_T_37) begin
      if (_T_11) begin
        out_ready_R_9 <= io_Out_9_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_9 <= 1'h0;
      end else if (_T_11) begin
        out_ready_R_9 <= io_Out_9_ready;
      end
    end else if (_T_11) begin
      out_ready_R_9 <= io_Out_9_ready;
    end
    if (reset) begin
      out_ready_R_10 <= 1'h0;
    end else if (_T_37) begin
      if (_T_12) begin
        out_ready_R_10 <= io_Out_10_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_10 <= 1'h0;
      end else if (_T_12) begin
        out_ready_R_10 <= io_Out_10_ready;
      end
    end else if (_T_12) begin
      out_ready_R_10 <= io_Out_10_ready;
    end
    if (reset) begin
      out_ready_R_11 <= 1'h0;
    end else if (_T_37) begin
      if (_T_13) begin
        out_ready_R_11 <= io_Out_11_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_11 <= 1'h0;
      end else if (_T_13) begin
        out_ready_R_11 <= io_Out_11_ready;
      end
    end else if (_T_13) begin
      out_ready_R_11 <= io_Out_11_ready;
    end
    if (reset) begin
      out_ready_R_12 <= 1'h0;
    end else if (_T_37) begin
      if (_T_14) begin
        out_ready_R_12 <= io_Out_12_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_12 <= 1'h0;
      end else if (_T_14) begin
        out_ready_R_12 <= io_Out_12_ready;
      end
    end else if (_T_14) begin
      out_ready_R_12 <= io_Out_12_ready;
    end
    if (reset) begin
      out_ready_R_13 <= 1'h0;
    end else if (_T_37) begin
      if (_T_15) begin
        out_ready_R_13 <= io_Out_13_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_13 <= 1'h0;
      end else if (_T_15) begin
        out_ready_R_13 <= io_Out_13_ready;
      end
    end else if (_T_15) begin
      out_ready_R_13 <= io_Out_13_ready;
    end
    if (reset) begin
      out_ready_R_14 <= 1'h0;
    end else if (_T_37) begin
      if (_T_16) begin
        out_ready_R_14 <= io_Out_14_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_14 <= 1'h0;
      end else if (_T_16) begin
        out_ready_R_14 <= io_Out_14_ready;
      end
    end else if (_T_16) begin
      out_ready_R_14 <= io_Out_14_ready;
    end
    if (reset) begin
      out_ready_R_15 <= 1'h0;
    end else if (_T_37) begin
      if (_T_17) begin
        out_ready_R_15 <= io_Out_15_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_15 <= 1'h0;
      end else if (_T_17) begin
        out_ready_R_15 <= io_Out_15_ready;
      end
    end else if (_T_17) begin
      out_ready_R_15 <= io_Out_15_ready;
    end
    if (reset) begin
      out_ready_R_16 <= 1'h0;
    end else if (_T_37) begin
      if (_T_18) begin
        out_ready_R_16 <= io_Out_16_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_16 <= 1'h0;
      end else if (_T_18) begin
        out_ready_R_16 <= io_Out_16_ready;
      end
    end else if (_T_18) begin
      out_ready_R_16 <= io_Out_16_ready;
    end
    if (reset) begin
      out_ready_R_17 <= 1'h0;
    end else if (_T_37) begin
      if (_T_19) begin
        out_ready_R_17 <= io_Out_17_ready;
      end
    end else if (state) begin
      if (_T_57) begin
        out_ready_R_17 <= 1'h0;
      end else if (_T_19) begin
        out_ready_R_17 <= io_Out_17_ready;
      end
    end else if (_T_19) begin
      out_ready_R_17 <= io_Out_17_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_0 <= _GEN_50;
    end else if (_T_2) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_1 <= _GEN_51;
    end else if (_T_3) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_2 <= _GEN_52;
    end else if (_T_4) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_3 <= _GEN_53;
    end else if (_T_5) begin
      out_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_4 <= _GEN_54;
    end else if (_T_6) begin
      out_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_5 <= _GEN_55;
    end else if (_T_7) begin
      out_valid_R_5 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_6 <= _GEN_56;
    end else if (_T_8) begin
      out_valid_R_6 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_7 <= _GEN_57;
    end else if (_T_9) begin
      out_valid_R_7 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_8 <= _GEN_58;
    end else if (_T_10) begin
      out_valid_R_8 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_9 <= _GEN_59;
    end else if (_T_11) begin
      out_valid_R_9 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_10 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_10 <= _GEN_60;
    end else if (_T_12) begin
      out_valid_R_10 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_11 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_11 <= _GEN_61;
    end else if (_T_13) begin
      out_valid_R_11 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_12 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_12 <= _GEN_62;
    end else if (_T_14) begin
      out_valid_R_12 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_13 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_13 <= _GEN_63;
    end else if (_T_15) begin
      out_valid_R_13 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_14 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_14 <= _GEN_64;
    end else if (_T_16) begin
      out_valid_R_14 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_15 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_15 <= _GEN_65;
    end else if (_T_17) begin
      out_valid_R_15 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_16 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_16 <= _GEN_66;
    end else if (_T_18) begin
      out_valid_R_16 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_17 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_17 <= _GEN_67;
    end else if (_T_19) begin
      out_valid_R_17 <= 1'h0;
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      mask_valid_R_0 <= _GEN_68;
    end else if (_T_20) begin
      mask_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_24;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else if (_T_28) begin
      predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else if (_T_28) begin
      predicate_in_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else if (_T_29) begin
      predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else if (_T_29) begin
      predicate_in_R_1_control <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else if (_T_28) begin
      predicate_control_R_0 <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else if (_T_29) begin
      predicate_control_R_1 <= io_predicateIn_1_bits_control;
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      predicate_valid_R_0 <= _T_30;
    end else if (state) begin
      if (_T_57) begin
        predicate_valid_R_0 <= 1'h0;
      end else begin
        predicate_valid_R_0 <= _T_30;
      end
    end else begin
      predicate_valid_R_0 <= _T_30;
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else if (_T_37) begin
      predicate_valid_R_1 <= _T_31;
    end else if (state) begin
      if (_T_57) begin
        predicate_valid_R_1 <= 1'h0;
      end else begin
        predicate_valid_R_1 <= _T_31;
      end
    end else begin
      predicate_valid_R_1 <= _T_31;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_37) begin
      state <= _GEN_69;
    end else if (state) begin
      if (_T_57) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_158 & _T_61) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] bb_for_body165] [Mask: 0x%x]\n",predicate_task,_T_36); // @[BasicBlock.scala 129:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_163 & _T_61) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] bb_for_body165: Output fired @ %d -> 0 predicate\n",cycleCount); // @[BasicBlock.scala 134:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_1(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 224:46]
  reg  in_data_R_0_control; // @[BasicBlock.scala 224:46]
  reg  in_data_valid_R_0; // @[BasicBlock.scala 225:52]
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 227:25]
  reg  output_valid_R_0; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_1; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_2; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_3; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_4; // @[BasicBlock.scala 228:49]
  reg  output_fire_R_0; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_1; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_2; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_3; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_4; // @[BasicBlock.scala 229:48]
  wire  _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 234:36]
  wire  _GEN_5 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 234:36]
  wire [4:0] in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 241:34]
  wire  _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 246:28]
  wire  _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 246:28]
  wire  _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_10 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 246:28]
  wire  _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 246:28]
  wire  _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 246:28]
  wire  out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 258:85]
  reg  state; // @[BasicBlock.scala 289:22]
  wire  _T_27 = ~state; // @[Conditional.scala 37:30]
  wire  _T_33 = _T_8 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_34 = _T_9 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_35 = _T_10 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_36 = _T_11 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_37 = _T_12 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_39 = ~reset; // @[BasicBlock.scala 311:17]
  wire  _GEN_16 = _GEN_5 | output_valid_R_0; // @[BasicBlock.scala 301:9]
  wire  _GEN_17 = _GEN_5 | output_valid_R_1; // @[BasicBlock.scala 301:9]
  wire  _GEN_18 = _GEN_5 | output_valid_R_2; // @[BasicBlock.scala 301:9]
  wire  _GEN_19 = _GEN_5 | output_valid_R_3; // @[BasicBlock.scala 301:9]
  wire  _GEN_20 = _GEN_5 | output_valid_R_4; // @[BasicBlock.scala 301:9]
  wire  _GEN_26 = _GEN_5 | state; // @[BasicBlock.scala 301:9]
  wire  _T_41 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 317:35]
  wire  _T_42 = _T_41 & out_fire_mask_2; // @[BasicBlock.scala 317:35]
  wire  _T_43 = _T_42 & out_fire_mask_3; // @[BasicBlock.scala 317:35]
  wire  _T_44 = _T_43 & out_fire_mask_4; // @[BasicBlock.scala 317:35]
  wire  _GEN_67 = _T_27 & _GEN_5; // @[BasicBlock.scala 311:17]
  assign io_predicateIn_0_ready = ~in_data_valid_R_0; // @[BasicBlock.scala 233:29]
  assign io_Out_0_valid = _T_27 ? _GEN_16 : output_valid_R_0; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_1_valid = _T_27 ? _GEN_17 : output_valid_R_1; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_2_valid = _T_27 ? _GEN_18 : output_valid_R_2; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_3_valid = _T_27 ? _GEN_19 : output_valid_R_3; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_4_valid = _T_27 ? _GEN_20 : output_valid_R_4; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_4_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (_T_7) begin
      in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_control <= 1'h0;
      end else if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (_T_7) begin
      in_data_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      in_data_valid_R_0 <= _GEN_5;
    end else if (state) begin
      if (_T_44) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_5;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_5;
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_0 <= _T_33;
      end else if (_T_8) begin
        output_valid_R_0 <= 1'h0;
      end
    end else if (_T_8) begin
      output_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_1 <= _T_34;
      end else if (_T_9) begin
        output_valid_R_1 <= 1'h0;
      end
    end else if (_T_9) begin
      output_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_2 <= _T_35;
      end else if (_T_10) begin
        output_valid_R_2 <= 1'h0;
      end
    end else if (_T_10) begin
      output_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_3 <= _T_36;
      end else if (_T_11) begin
        output_valid_R_3 <= 1'h0;
      end
    end else if (_T_11) begin
      output_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_4 <= _T_37;
      end else if (_T_12) begin
        output_valid_R_4 <= 1'h0;
      end
    end else if (_T_12) begin
      output_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_0 <= _GEN_6;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_0 <= 1'h0;
      end else begin
        output_fire_R_0 <= _GEN_6;
      end
    end else begin
      output_fire_R_0 <= _GEN_6;
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_1 <= _GEN_8;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_1 <= 1'h0;
      end else begin
        output_fire_R_1 <= _GEN_8;
      end
    end else begin
      output_fire_R_1 <= _GEN_8;
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_2 <= _GEN_10;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_2 <= 1'h0;
      end else begin
        output_fire_R_2 <= _GEN_10;
      end
    end else begin
      output_fire_R_2 <= _GEN_10;
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_3 <= _GEN_12;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_3 <= 1'h0;
      end else begin
        output_fire_R_3 <= _GEN_12;
      end
    end else begin
      output_fire_R_3 <= _GEN_12;
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_4 <= _GEN_14;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_4 <= 1'h0;
      end else begin
        output_fire_R_4 <= _GEN_14;
      end
    end else begin
      output_fire_R_4 <= _GEN_14;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_27) begin
      state <= _GEN_26;
    end else if (state) begin
      if (_T_44) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] [bb_for_inc276] [Out: %d] [Cycle: %d]\n",output_R_taskID,_GEN_3,cycleCount); // @[BasicBlock.scala 311:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_2(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 224:46]
  reg  in_data_R_0_control; // @[BasicBlock.scala 224:46]
  reg  in_data_valid_R_0; // @[BasicBlock.scala 225:52]
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 227:25]
  reg  output_valid_R_0; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_1; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_2; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_3; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_4; // @[BasicBlock.scala 228:49]
  reg  output_fire_R_0; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_1; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_2; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_3; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_4; // @[BasicBlock.scala 229:48]
  wire  _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 234:36]
  wire  _GEN_5 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 234:36]
  wire [4:0] in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 241:34]
  wire  _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 246:28]
  wire  _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 246:28]
  wire  _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_10 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 246:28]
  wire  _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 246:28]
  wire  _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 246:28]
  wire  out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 258:85]
  reg  state; // @[BasicBlock.scala 289:22]
  wire  _T_27 = ~state; // @[Conditional.scala 37:30]
  wire  _T_33 = _T_8 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_34 = _T_9 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_35 = _T_10 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_36 = _T_11 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_37 = _T_12 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_39 = ~reset; // @[BasicBlock.scala 311:17]
  wire  _GEN_16 = _GEN_5 | output_valid_R_0; // @[BasicBlock.scala 301:9]
  wire  _GEN_17 = _GEN_5 | output_valid_R_1; // @[BasicBlock.scala 301:9]
  wire  _GEN_18 = _GEN_5 | output_valid_R_2; // @[BasicBlock.scala 301:9]
  wire  _GEN_19 = _GEN_5 | output_valid_R_3; // @[BasicBlock.scala 301:9]
  wire  _GEN_20 = _GEN_5 | output_valid_R_4; // @[BasicBlock.scala 301:9]
  wire  _GEN_26 = _GEN_5 | state; // @[BasicBlock.scala 301:9]
  wire  _T_41 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 317:35]
  wire  _T_42 = _T_41 & out_fire_mask_2; // @[BasicBlock.scala 317:35]
  wire  _T_43 = _T_42 & out_fire_mask_3; // @[BasicBlock.scala 317:35]
  wire  _T_44 = _T_43 & out_fire_mask_4; // @[BasicBlock.scala 317:35]
  wire  _GEN_67 = _T_27 & _GEN_5; // @[BasicBlock.scala 311:17]
  assign io_predicateIn_0_ready = ~in_data_valid_R_0; // @[BasicBlock.scala 233:29]
  assign io_Out_0_valid = _T_27 ? _GEN_16 : output_valid_R_0; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_1_valid = _T_27 ? _GEN_17 : output_valid_R_1; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_2_valid = _T_27 ? _GEN_18 : output_valid_R_2; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_3_valid = _T_27 ? _GEN_19 : output_valid_R_3; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_4_valid = _T_27 ? _GEN_20 : output_valid_R_4; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_4_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (_T_7) begin
      in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_control <= 1'h0;
      end else if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (_T_7) begin
      in_data_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      in_data_valid_R_0 <= _GEN_5;
    end else if (state) begin
      if (_T_44) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_5;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_5;
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_0 <= _T_33;
      end else if (_T_8) begin
        output_valid_R_0 <= 1'h0;
      end
    end else if (_T_8) begin
      output_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_1 <= _T_34;
      end else if (_T_9) begin
        output_valid_R_1 <= 1'h0;
      end
    end else if (_T_9) begin
      output_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_2 <= _T_35;
      end else if (_T_10) begin
        output_valid_R_2 <= 1'h0;
      end
    end else if (_T_10) begin
      output_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_3 <= _T_36;
      end else if (_T_11) begin
        output_valid_R_3 <= 1'h0;
      end
    end else if (_T_11) begin
      output_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_4 <= _T_37;
      end else if (_T_12) begin
        output_valid_R_4 <= 1'h0;
      end
    end else if (_T_12) begin
      output_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_0 <= _GEN_6;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_0 <= 1'h0;
      end else begin
        output_fire_R_0 <= _GEN_6;
      end
    end else begin
      output_fire_R_0 <= _GEN_6;
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_1 <= _GEN_8;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_1 <= 1'h0;
      end else begin
        output_fire_R_1 <= _GEN_8;
      end
    end else begin
      output_fire_R_1 <= _GEN_8;
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_2 <= _GEN_10;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_2 <= 1'h0;
      end else begin
        output_fire_R_2 <= _GEN_10;
      end
    end else begin
      output_fire_R_2 <= _GEN_10;
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_3 <= _GEN_12;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_3 <= 1'h0;
      end else begin
        output_fire_R_3 <= _GEN_12;
      end
    end else begin
      output_fire_R_3 <= _GEN_12;
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_4 <= _GEN_14;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_4 <= 1'h0;
      end else begin
        output_fire_R_4 <= _GEN_14;
      end
    end else begin
      output_fire_R_4 <= _GEN_14;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_27) begin
      state <= _GEN_26;
    end else if (state) begin
      if (_T_44) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] [bb_for_inc307] [Out: %d] [Cycle: %d]\n",output_R_taskID,_GEN_3,cycleCount); // @[BasicBlock.scala 311:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_3(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 224:46]
  reg  in_data_R_0_control; // @[BasicBlock.scala 224:46]
  reg  in_data_valid_R_0; // @[BasicBlock.scala 225:52]
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 227:25]
  reg  output_valid_R_0; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_1; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_2; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_3; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_4; // @[BasicBlock.scala 228:49]
  reg  output_fire_R_0; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_1; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_2; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_3; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_4; // @[BasicBlock.scala 229:48]
  wire  _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 234:36]
  wire  _GEN_5 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 234:36]
  wire [4:0] in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 241:34]
  wire  _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 246:28]
  wire  _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 246:28]
  wire  _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_10 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 246:28]
  wire  _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 246:28]
  wire  _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 246:28]
  wire  out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 258:85]
  reg  state; // @[BasicBlock.scala 289:22]
  wire  _T_27 = ~state; // @[Conditional.scala 37:30]
  wire  _T_33 = _T_8 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_34 = _T_9 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_35 = _T_10 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_36 = _T_11 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_37 = _T_12 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_39 = ~reset; // @[BasicBlock.scala 311:17]
  wire  _GEN_16 = _GEN_5 | output_valid_R_0; // @[BasicBlock.scala 301:9]
  wire  _GEN_17 = _GEN_5 | output_valid_R_1; // @[BasicBlock.scala 301:9]
  wire  _GEN_18 = _GEN_5 | output_valid_R_2; // @[BasicBlock.scala 301:9]
  wire  _GEN_19 = _GEN_5 | output_valid_R_3; // @[BasicBlock.scala 301:9]
  wire  _GEN_20 = _GEN_5 | output_valid_R_4; // @[BasicBlock.scala 301:9]
  wire  _GEN_26 = _GEN_5 | state; // @[BasicBlock.scala 301:9]
  wire  _T_41 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 317:35]
  wire  _T_42 = _T_41 & out_fire_mask_2; // @[BasicBlock.scala 317:35]
  wire  _T_43 = _T_42 & out_fire_mask_3; // @[BasicBlock.scala 317:35]
  wire  _T_44 = _T_43 & out_fire_mask_4; // @[BasicBlock.scala 317:35]
  wire  _GEN_67 = _T_27 & _GEN_5; // @[BasicBlock.scala 311:17]
  assign io_predicateIn_0_ready = ~in_data_valid_R_0; // @[BasicBlock.scala 233:29]
  assign io_Out_0_valid = _T_27 ? _GEN_16 : output_valid_R_0; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_1_valid = _T_27 ? _GEN_17 : output_valid_R_1; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_2_valid = _T_27 ? _GEN_18 : output_valid_R_2; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_3_valid = _T_27 ? _GEN_19 : output_valid_R_3; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_4_valid = _T_27 ? _GEN_20 : output_valid_R_4; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_4_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (_T_7) begin
      in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_control <= 1'h0;
      end else if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (_T_7) begin
      in_data_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      in_data_valid_R_0 <= _GEN_5;
    end else if (state) begin
      if (_T_44) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_5;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_5;
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_0 <= _T_33;
      end else if (_T_8) begin
        output_valid_R_0 <= 1'h0;
      end
    end else if (_T_8) begin
      output_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_1 <= _T_34;
      end else if (_T_9) begin
        output_valid_R_1 <= 1'h0;
      end
    end else if (_T_9) begin
      output_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_2 <= _T_35;
      end else if (_T_10) begin
        output_valid_R_2 <= 1'h0;
      end
    end else if (_T_10) begin
      output_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_3 <= _T_36;
      end else if (_T_11) begin
        output_valid_R_3 <= 1'h0;
      end
    end else if (_T_11) begin
      output_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_4 <= _T_37;
      end else if (_T_12) begin
        output_valid_R_4 <= 1'h0;
      end
    end else if (_T_12) begin
      output_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_0 <= _GEN_6;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_0 <= 1'h0;
      end else begin
        output_fire_R_0 <= _GEN_6;
      end
    end else begin
      output_fire_R_0 <= _GEN_6;
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_1 <= _GEN_8;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_1 <= 1'h0;
      end else begin
        output_fire_R_1 <= _GEN_8;
      end
    end else begin
      output_fire_R_1 <= _GEN_8;
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_2 <= _GEN_10;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_2 <= 1'h0;
      end else begin
        output_fire_R_2 <= _GEN_10;
      end
    end else begin
      output_fire_R_2 <= _GEN_10;
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_3 <= _GEN_12;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_3 <= 1'h0;
      end else begin
        output_fire_R_3 <= _GEN_12;
      end
    end else begin
      output_fire_R_3 <= _GEN_12;
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_4 <= _GEN_14;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_4 <= 1'h0;
      end else begin
        output_fire_R_4 <= _GEN_14;
      end
    end else begin
      output_fire_R_4 <= _GEN_14;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_27) begin
      state <= _GEN_26;
    end else if (state) begin
      if (_T_44) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] [bb_for_inc338] [Out: %d] [Cycle: %d]\n",output_R_taskID,_GEN_3,cycleCount); // @[BasicBlock.scala 311:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_4(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 224:46]
  reg  in_data_R_0_control; // @[BasicBlock.scala 224:46]
  reg  in_data_valid_R_0; // @[BasicBlock.scala 225:52]
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 227:25]
  reg  output_valid_R_0; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_1; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_2; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_3; // @[BasicBlock.scala 228:49]
  reg  output_valid_R_4; // @[BasicBlock.scala 228:49]
  reg  output_fire_R_0; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_1; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_2; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_3; // @[BasicBlock.scala 229:48]
  reg  output_fire_R_4; // @[BasicBlock.scala 229:48]
  wire  _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 234:36]
  wire  _GEN_5 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 234:36]
  wire [4:0] in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 241:34]
  wire  _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 246:28]
  wire  _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 246:28]
  wire  _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_10 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 246:28]
  wire  _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 246:28]
  wire  _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 246:28]
  wire  out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 258:85]
  wire  out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 258:85]
  reg  state; // @[BasicBlock.scala 289:22]
  wire  _T_27 = ~state; // @[Conditional.scala 37:30]
  wire  _T_33 = _T_8 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_34 = _T_9 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_35 = _T_10 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_36 = _T_11 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_37 = _T_12 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_39 = ~reset; // @[BasicBlock.scala 311:17]
  wire  _GEN_16 = _GEN_5 | output_valid_R_0; // @[BasicBlock.scala 301:9]
  wire  _GEN_17 = _GEN_5 | output_valid_R_1; // @[BasicBlock.scala 301:9]
  wire  _GEN_18 = _GEN_5 | output_valid_R_2; // @[BasicBlock.scala 301:9]
  wire  _GEN_19 = _GEN_5 | output_valid_R_3; // @[BasicBlock.scala 301:9]
  wire  _GEN_20 = _GEN_5 | output_valid_R_4; // @[BasicBlock.scala 301:9]
  wire  _GEN_26 = _GEN_5 | state; // @[BasicBlock.scala 301:9]
  wire  _T_41 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 317:35]
  wire  _T_42 = _T_41 & out_fire_mask_2; // @[BasicBlock.scala 317:35]
  wire  _T_43 = _T_42 & out_fire_mask_3; // @[BasicBlock.scala 317:35]
  wire  _T_44 = _T_43 & out_fire_mask_4; // @[BasicBlock.scala 317:35]
  wire  _GEN_67 = _T_27 & _GEN_5; // @[BasicBlock.scala 311:17]
  assign io_predicateIn_0_ready = ~in_data_valid_R_0; // @[BasicBlock.scala 233:29]
  assign io_Out_0_valid = _T_27 ? _GEN_16 : output_valid_R_0; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_1_valid = _T_27 ? _GEN_17 : output_valid_R_1; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_2_valid = _T_27 ? _GEN_18 : output_valid_R_2; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_3_valid = _T_27 ? _GEN_19 : output_valid_R_3; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
  assign io_Out_4_valid = _T_27 ? _GEN_20 : output_valid_R_4; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
  assign io_Out_4_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 279:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (_T_7) begin
      in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else if (_T_27) begin
      if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (state) begin
      if (_T_44) begin
        in_data_R_0_control <= 1'h0;
      end else if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (_T_7) begin
      in_data_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      in_data_valid_R_0 <= _GEN_5;
    end else if (state) begin
      if (_T_44) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_5;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_5;
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_0 <= _T_33;
      end else if (_T_8) begin
        output_valid_R_0 <= 1'h0;
      end
    end else if (_T_8) begin
      output_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_1 <= _T_34;
      end else if (_T_9) begin
        output_valid_R_1 <= 1'h0;
      end
    end else if (_T_9) begin
      output_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_2 <= _T_35;
      end else if (_T_10) begin
        output_valid_R_2 <= 1'h0;
      end
    end else if (_T_10) begin
      output_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_3 <= _T_36;
      end else if (_T_11) begin
        output_valid_R_3 <= 1'h0;
      end
    end else if (_T_11) begin
      output_valid_R_3 <= 1'h0;
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else if (_T_27) begin
      if (_GEN_5) begin
        output_valid_R_4 <= _T_37;
      end else if (_T_12) begin
        output_valid_R_4 <= 1'h0;
      end
    end else if (_T_12) begin
      output_valid_R_4 <= 1'h0;
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_0 <= _GEN_6;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_0 <= 1'h0;
      end else begin
        output_fire_R_0 <= _GEN_6;
      end
    end else begin
      output_fire_R_0 <= _GEN_6;
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_1 <= _GEN_8;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_1 <= 1'h0;
      end else begin
        output_fire_R_1 <= _GEN_8;
      end
    end else begin
      output_fire_R_1 <= _GEN_8;
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_2 <= _GEN_10;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_2 <= 1'h0;
      end else begin
        output_fire_R_2 <= _GEN_10;
      end
    end else begin
      output_fire_R_2 <= _GEN_10;
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_3 <= _GEN_12;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_3 <= 1'h0;
      end else begin
        output_fire_R_3 <= _GEN_12;
      end
    end else begin
      output_fire_R_3 <= _GEN_12;
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else if (_T_27) begin
      output_fire_R_4 <= _GEN_14;
    end else if (state) begin
      if (_T_44) begin
        output_fire_R_4 <= 1'h0;
      end else begin
        output_fire_R_4 <= _GEN_14;
      end
    end else begin
      output_fire_R_4 <= _GEN_14;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_27) begin
      state <= _GEN_26;
    end else if (state) begin
      if (_T_44) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] [bb_for_inc369] [Out: %d] [Cycle: %d]\n",output_R_taskID,_GEN_3,cycleCount); // @[BasicBlock.scala 311:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_5(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 224:46]
  reg  in_data_R_0_control; // @[BasicBlock.scala 224:46]
  reg  in_data_valid_R_0; // @[BasicBlock.scala 225:52]
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 227:25]
  reg  output_valid_R_0; // @[BasicBlock.scala 228:49]
  reg  output_fire_R_0; // @[BasicBlock.scala 229:48]
  wire  _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 234:36]
  wire  _GEN_5 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 234:36]
  wire [4:0] in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 241:34]
  wire  _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_6 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 246:28]
  wire  out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 258:85]
  reg  state; // @[BasicBlock.scala 289:22]
  wire  _T_15 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 306:81]
  wire  _T_19 = ~reset; // @[BasicBlock.scala 311:17]
  wire  _GEN_8 = _GEN_5 | output_valid_R_0; // @[BasicBlock.scala 301:9]
  wire  _GEN_10 = _GEN_5 | state; // @[BasicBlock.scala 301:9]
  wire  _GEN_31 = _T_15 & _GEN_5; // @[BasicBlock.scala 311:17]
  assign io_predicateIn_0_ready = ~in_data_valid_R_0; // @[BasicBlock.scala 233:29]
  assign io_Out_0_valid = _T_15 ? _GEN_8 : output_valid_R_0; // @[BasicBlock.scala 284:21 BasicBlock.scala 303:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 279:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_15) begin
      if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (state) begin
      if (out_fire_mask_0) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_7) begin
        in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end else if (_T_7) begin
      in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else if (_T_15) begin
      if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (state) begin
      if (out_fire_mask_0) begin
        in_data_R_0_control <= 1'h0;
      end else if (_T_7) begin
        in_data_R_0_control <= io_predicateIn_0_bits_control;
      end
    end else if (_T_7) begin
      in_data_R_0_control <= io_predicateIn_0_bits_control;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      in_data_valid_R_0 <= _GEN_5;
    end else if (state) begin
      if (out_fire_mask_0) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_5;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_5;
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      if (_GEN_5) begin
        output_valid_R_0 <= _T_17;
      end else if (_T_8) begin
        output_valid_R_0 <= 1'h0;
      end
    end else if (_T_8) begin
      output_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else if (_T_15) begin
      output_fire_R_0 <= _GEN_6;
    end else if (state) begin
      if (out_fire_mask_0) begin
        output_fire_R_0 <= 1'h0;
      end else begin
        output_fire_R_0 <= _GEN_6;
      end
    end else begin
      output_fire_R_0 <= _GEN_6;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_15) begin
      state <= _GEN_10;
    end else if (state) begin
      if (out_fire_mask_0) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [BB] [bb_for_end3810] [Out: %d] [Cycle: %d]\n",output_R_taskID,_GEN_3,cycleCount); // @[BasicBlock.scala 311:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode(
  input   clock,
  input   reset,
  output  io_enable_ready,
  input   io_enable_valid,
  input   io_enable_bits_control,
  input   io_Out_0_ready,
  output  io_Out_0_valid,
  output  io_Out_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  state; // @[BranchNode.scala 588:22]
  wire  _T_11 = ~state; // @[Conditional.scala 37:30]
  wire  _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_16 = ~reset; // @[BranchNode.scala 616:17]
  wire  _GEN_8 = enable_valid_R | state; // @[BranchNode.scala 611:46]
  wire  _GEN_10 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 611:46]
  wire  _T_18 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_19 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_20 = _T_18 | _T_19; // @[HandShaking.scala 725:29]
  wire  _GEN_31 = _T_11 & enable_valid_R; // @[BranchNode.scala 616:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = _T_11 ? _GEN_10 : out_valid_R_0; // @[HandShaking.scala 630:21 BranchNode.scala 614:32]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 607:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cycleCount = _RAND_4[14:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_control <= 1'h0;
      end else if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_20) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (enable_valid_R) begin
        out_valid_R_0 <= _T_14;
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_11) begin
      state <= _GEN_8;
    end else if (state) begin
      if (_T_20) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [UBR] [br_0] [Out: %d] [Cycle: %d]\n",5'h0,enable_R_control,cycleCount); // @[BranchNode.scala 616:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [63:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[PhiNode.scala 203:26]
  reg [4:0] in_data_R_1_taskID; // @[PhiNode.scala 203:26]
  reg [63:0] in_data_R_1_data; // @[PhiNode.scala 203:26]
  reg  in_data_valid_R_0; // @[PhiNode.scala 204:32]
  reg  in_data_valid_R_1; // @[PhiNode.scala 204:32]
  reg  enable_R_control; // @[PhiNode.scala 207:25]
  reg  enable_valid_R; // @[PhiNode.scala 208:31]
  reg [1:0] mask_R; // @[PhiNode.scala 211:23]
  reg  mask_valid_R; // @[PhiNode.scala 212:29]
  reg [1:0] state; // @[PhiNode.scala 216:22]
  reg  out_valid_R_0; // @[PhiNode.scala 219:49]
  reg  out_valid_R_1; // @[PhiNode.scala 219:49]
  reg  fire_R_0; // @[PhiNode.scala 221:44]
  reg  fire_R_1; // @[PhiNode.scala 221:44]
  wire  _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_10 | mask_valid_R; // @[PhiNode.scala 239:24]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_12 | enable_valid_R; // @[PhiNode.scala 246:26]
  wire  _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 254:29]
  wire  _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 254:29]
  wire  sel = mask_R[1]; // @[CircuitMath.scala 30:8]
  wire  _T_17 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_16 = _T_17 | fire_R_0; // @[PhiNode.scala 276:26]
  wire  _GEN_17 = _T_17 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 276:26]
  wire  _T_18 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = _T_18 | fire_R_1; // @[PhiNode.scala 276:26]
  wire  _GEN_19 = _T_18 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 276:26]
  wire  fire_mask_0 = fire_R_0 | _T_17; // @[PhiNode.scala 283:74]
  wire  fire_mask_1 = fire_R_1 | _T_18; // @[PhiNode.scala 283:74]
  wire [63:0] _GEN_27 = sel ? in_data_R_1_data : 64'h0; // @[PhiNode.scala 312:12]
  wire  _T_38 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_39 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 286:30]
  wire  _T_40 = enable_valid_R & _T_39; // @[PhiNode.scala 327:27]
  reg [2:0] guard_index; // @[Counter.scala 29:33]
  wire [63:0] _GEN_29 = 3'h1 == guard_index ? 64'h2 : 64'h0; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_30 = 3'h2 == guard_index ? 64'h4 : _GEN_29; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_31 = 3'h3 == guard_index ? 64'h6 : _GEN_30; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_32 = 3'h4 == guard_index ? 64'h8 : _GEN_31; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_33 = 3'h5 == guard_index ? 64'ha : _GEN_32; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_34 = 3'h6 == guard_index ? 64'hc : _GEN_33; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_35 = 3'h7 == guard_index ? 64'he : _GEN_34; // @[PhiNode.scala 336:38]
  wire  _T_42 = _GEN_27 != _GEN_35; // @[PhiNode.scala 336:38]
  wire  _T_31 = _T_40 & enable_R_control; // @[PhiNode.scala 290:38]
  wire  _T_32 = state == 2'h0; // @[PhiNode.scala 290:67]
  wire  _T_33 = _T_31 & _T_32; // @[PhiNode.scala 290:58]
  wire [2:0] _T_37 = guard_index + 3'h1; // @[Counter.scala 39:22]
  wire [4:0] _GEN_26 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 312:12]
  wire  _T_44 = ~reset; // @[PhiNode.scala 341:23]
  wire [4:0] _GEN_46 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 350:19]
  wire  _GEN_51 = _T_40 | _GEN_17; // @[PhiNode.scala 327:66]
  wire  _GEN_52 = _T_40 | _GEN_19; // @[PhiNode.scala 327:66]
  wire  _T_49 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_50 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 364:31]
  wire  _T_54 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_91 = _T_54 ? 64'h0 : _GEN_27; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_132 = _T_49 ? _GEN_27 : _GEN_91; // @[Conditional.scala 39:67]
  wire  _GEN_165 = _T_38 & _T_40; // @[PhiNode.scala 341:23]
  wire  _GEN_166 = _GEN_165 & enable_R_control; // @[PhiNode.scala 341:23]
  wire  _GEN_167 = _GEN_166 & _T_42; // @[PhiNode.scala 341:23]
  wire  _GEN_171 = ~enable_R_control; // @[PhiNode.scala 357:19]
  wire  _GEN_172 = _GEN_165 & _GEN_171; // @[PhiNode.scala 357:19]
  assign io_enable_ready = ~enable_valid_R; // @[PhiNode.scala 245:19]
  assign io_InData_0_ready = ~in_data_valid_R_0; // @[PhiNode.scala 253:24]
  assign io_InData_1_ready = ~in_data_valid_R_1; // @[PhiNode.scala 253:24]
  assign io_Mask_ready = ~mask_valid_R; // @[PhiNode.scala 238:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 322:21]
  assign io_Out_0_bits_data = _T_38 ? _GEN_27 : _GEN_132; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 322:21]
  assign io_Out_1_bits_data = _T_38 ? _GEN_27 : _GEN_132; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[4:0];
  _RAND_3 = {2{`RANDOM}};
  in_data_R_1_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_R_control = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enable_valid_R = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mask_R = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  mask_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fire_R_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  guard_index = _RAND_15[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_14) begin
      in_data_R_0_taskID <= io_InData_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_R_1_taskID <= 5'h0;
      end else if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_R_1_taskID <= 5'h0;
      end else if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_16) begin
      in_data_R_1_taskID <= io_InData_1_bits_taskID;
    end
    if (reset) begin
      in_data_R_1_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_16) begin
      in_data_R_1_data <= io_InData_1_bits_data;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      in_data_valid_R_0 <= _GEN_11;
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_11;
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else if (_T_38) begin
      in_data_valid_R_1 <= _GEN_15;
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else begin
      in_data_valid_R_1 <= _GEN_15;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_38) begin
      enable_valid_R <= _GEN_7;
    end else if (_T_49) begin
      if (_T_50) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else begin
      enable_valid_R <= _GEN_7;
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else if (_T_38) begin
      if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_10) begin
      mask_R <= io_Mask_bits;
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else if (_T_38) begin
      mask_valid_R <= _GEN_3;
    end else if (_T_49) begin
      if (_T_50) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else begin
      mask_valid_R <= _GEN_3;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_38) begin
      if (_T_40) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_49) begin
      if (_T_50) begin
        state <= 2'h0;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      out_valid_R_0 <= _GEN_51;
    end else if (_T_17) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_38) begin
      out_valid_R_1 <= _GEN_52;
    end else if (_T_18) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else if (_T_38) begin
      fire_R_0 <= _GEN_16;
    end else if (_T_49) begin
      if (_T_50) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else begin
      fire_R_0 <= _GEN_16;
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else if (_T_38) begin
      fire_R_1 <= _GEN_18;
    end else if (_T_49) begin
      if (_T_50) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else begin
      fire_R_1 <= _GEN_18;
    end
    if (reset) begin
      guard_index <= 3'h0;
    end else if (_T_33) begin
      guard_index <= _T_37;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_167 & _T_44) begin
          $fwrite(32'h80000002,"[DEBUG] [Bbgemm] [TID->%d] [PHI] phiindvars_iv841 Produced value: %d, correct value: %d\n",_GEN_26,_GEN_27,_GEN_35); // @[PhiNode.scala 341:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_166 & _T_44) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv841] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_46,enable_R_control,_GEN_27,cycleCount); // @[PhiNode.scala 350:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_172 & _T_44) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv841] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_46,enable_R_control,_GEN_27,cycleCount); // @[PhiNode.scala 357:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_1(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  state; // @[BranchNode.scala 588:22]
  wire  _T_11 = ~state; // @[Conditional.scala 37:30]
  wire  _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_16 = ~reset; // @[BranchNode.scala 616:17]
  wire  _GEN_8 = enable_valid_R | state; // @[BranchNode.scala 611:46]
  wire  _GEN_10 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 611:46]
  wire  _T_18 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_19 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_20 = _T_18 | _T_19; // @[HandShaking.scala 725:29]
  wire  _GEN_31 = _T_11 & enable_valid_R; // @[BranchNode.scala 616:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = _T_11 ? _GEN_10 : out_valid_R_0; // @[HandShaking.scala 630:21 BranchNode.scala 614:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 607:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 607:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_control <= 1'h0;
      end else if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_20) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (enable_valid_R) begin
        out_valid_R_0 <= _T_14;
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_11) begin
      state <= _GEN_8;
    end else if (state) begin
      if (_T_20) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [UBR] [br_2] [Out: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,cycleCount); // @[BranchNode.scala 616:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [63:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[PhiNode.scala 203:26]
  reg [4:0] in_data_R_1_taskID; // @[PhiNode.scala 203:26]
  reg [63:0] in_data_R_1_data; // @[PhiNode.scala 203:26]
  reg  in_data_valid_R_0; // @[PhiNode.scala 204:32]
  reg  in_data_valid_R_1; // @[PhiNode.scala 204:32]
  reg  enable_R_control; // @[PhiNode.scala 207:25]
  reg  enable_valid_R; // @[PhiNode.scala 208:31]
  reg [1:0] mask_R; // @[PhiNode.scala 211:23]
  reg  mask_valid_R; // @[PhiNode.scala 212:29]
  reg [1:0] state; // @[PhiNode.scala 216:22]
  reg  out_valid_R_0; // @[PhiNode.scala 219:49]
  reg  out_valid_R_1; // @[PhiNode.scala 219:49]
  reg  fire_R_0; // @[PhiNode.scala 221:44]
  reg  fire_R_1; // @[PhiNode.scala 221:44]
  wire  _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_10 | mask_valid_R; // @[PhiNode.scala 239:24]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_12 | enable_valid_R; // @[PhiNode.scala 246:26]
  wire  _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 254:29]
  wire  _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 254:29]
  wire  sel = mask_R[1]; // @[CircuitMath.scala 30:8]
  wire  _T_17 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_16 = _T_17 | fire_R_0; // @[PhiNode.scala 276:26]
  wire  _GEN_17 = _T_17 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 276:26]
  wire  _T_18 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = _T_18 | fire_R_1; // @[PhiNode.scala 276:26]
  wire  _GEN_19 = _T_18 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 276:26]
  wire  fire_mask_0 = fire_R_0 | _T_17; // @[PhiNode.scala 283:74]
  wire  fire_mask_1 = fire_R_1 | _T_18; // @[PhiNode.scala 283:74]
  wire [63:0] _GEN_27 = sel ? in_data_R_1_data : 64'h0; // @[PhiNode.scala 312:12]
  wire  _T_38 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_39 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 286:30]
  wire  _T_40 = enable_valid_R & _T_39; // @[PhiNode.scala 327:27]
  reg [5:0] guard_index; // @[Counter.scala 29:33]
  wire [63:0] _GEN_29 = 6'h1 == guard_index ? 64'h2 : 64'h0; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_30 = 6'h2 == guard_index ? 64'h4 : _GEN_29; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_31 = 6'h3 == guard_index ? 64'h6 : _GEN_30; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_32 = 6'h4 == guard_index ? 64'h8 : _GEN_31; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_33 = 6'h5 == guard_index ? 64'ha : _GEN_32; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_34 = 6'h6 == guard_index ? 64'hc : _GEN_33; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_35 = 6'h7 == guard_index ? 64'he : _GEN_34; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_36 = 6'h8 == guard_index ? 64'h0 : _GEN_35; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_37 = 6'h9 == guard_index ? 64'h2 : _GEN_36; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_38 = 6'ha == guard_index ? 64'h4 : _GEN_37; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_39 = 6'hb == guard_index ? 64'h6 : _GEN_38; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_40 = 6'hc == guard_index ? 64'h8 : _GEN_39; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_41 = 6'hd == guard_index ? 64'ha : _GEN_40; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_42 = 6'he == guard_index ? 64'hc : _GEN_41; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_43 = 6'hf == guard_index ? 64'he : _GEN_42; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_44 = 6'h10 == guard_index ? 64'h0 : _GEN_43; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_45 = 6'h11 == guard_index ? 64'h2 : _GEN_44; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_46 = 6'h12 == guard_index ? 64'h4 : _GEN_45; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_47 = 6'h13 == guard_index ? 64'h6 : _GEN_46; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_48 = 6'h14 == guard_index ? 64'h8 : _GEN_47; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_49 = 6'h15 == guard_index ? 64'ha : _GEN_48; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_50 = 6'h16 == guard_index ? 64'hc : _GEN_49; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_51 = 6'h17 == guard_index ? 64'he : _GEN_50; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_52 = 6'h18 == guard_index ? 64'h0 : _GEN_51; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_53 = 6'h19 == guard_index ? 64'h2 : _GEN_52; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_54 = 6'h1a == guard_index ? 64'h4 : _GEN_53; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_55 = 6'h1b == guard_index ? 64'h6 : _GEN_54; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_56 = 6'h1c == guard_index ? 64'h8 : _GEN_55; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_57 = 6'h1d == guard_index ? 64'ha : _GEN_56; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_58 = 6'h1e == guard_index ? 64'hc : _GEN_57; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_59 = 6'h1f == guard_index ? 64'he : _GEN_58; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_60 = 6'h20 == guard_index ? 64'h0 : _GEN_59; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_61 = 6'h21 == guard_index ? 64'h2 : _GEN_60; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_62 = 6'h22 == guard_index ? 64'h4 : _GEN_61; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_63 = 6'h23 == guard_index ? 64'h6 : _GEN_62; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_64 = 6'h24 == guard_index ? 64'h8 : _GEN_63; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_65 = 6'h25 == guard_index ? 64'ha : _GEN_64; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_66 = 6'h26 == guard_index ? 64'hc : _GEN_65; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_67 = 6'h27 == guard_index ? 64'he : _GEN_66; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_68 = 6'h28 == guard_index ? 64'h0 : _GEN_67; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_69 = 6'h29 == guard_index ? 64'h2 : _GEN_68; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_70 = 6'h2a == guard_index ? 64'h4 : _GEN_69; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_71 = 6'h2b == guard_index ? 64'h6 : _GEN_70; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_72 = 6'h2c == guard_index ? 64'h8 : _GEN_71; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_73 = 6'h2d == guard_index ? 64'ha : _GEN_72; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_74 = 6'h2e == guard_index ? 64'hc : _GEN_73; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_75 = 6'h2f == guard_index ? 64'he : _GEN_74; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_76 = 6'h30 == guard_index ? 64'h0 : _GEN_75; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_77 = 6'h31 == guard_index ? 64'h2 : _GEN_76; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_78 = 6'h32 == guard_index ? 64'h4 : _GEN_77; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_79 = 6'h33 == guard_index ? 64'h6 : _GEN_78; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_80 = 6'h34 == guard_index ? 64'h8 : _GEN_79; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_81 = 6'h35 == guard_index ? 64'ha : _GEN_80; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_82 = 6'h36 == guard_index ? 64'hc : _GEN_81; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_83 = 6'h37 == guard_index ? 64'he : _GEN_82; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_84 = 6'h38 == guard_index ? 64'h0 : _GEN_83; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_85 = 6'h39 == guard_index ? 64'h2 : _GEN_84; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_86 = 6'h3a == guard_index ? 64'h4 : _GEN_85; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_87 = 6'h3b == guard_index ? 64'h6 : _GEN_86; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_88 = 6'h3c == guard_index ? 64'h8 : _GEN_87; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_89 = 6'h3d == guard_index ? 64'ha : _GEN_88; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_90 = 6'h3e == guard_index ? 64'hc : _GEN_89; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_91 = 6'h3f == guard_index ? 64'he : _GEN_90; // @[PhiNode.scala 336:38]
  wire  _T_42 = _GEN_27 != _GEN_91; // @[PhiNode.scala 336:38]
  wire  _T_31 = _T_40 & enable_R_control; // @[PhiNode.scala 290:38]
  wire  _T_32 = state == 2'h0; // @[PhiNode.scala 290:67]
  wire  _T_33 = _T_31 & _T_32; // @[PhiNode.scala 290:58]
  wire [5:0] _T_37 = guard_index + 6'h1; // @[Counter.scala 39:22]
  wire [4:0] _GEN_26 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 312:12]
  wire  _T_44 = ~reset; // @[PhiNode.scala 341:23]
  wire [4:0] _GEN_102 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 350:19]
  wire  _GEN_107 = _T_40 | _GEN_17; // @[PhiNode.scala 327:66]
  wire  _GEN_108 = _T_40 | _GEN_19; // @[PhiNode.scala 327:66]
  wire  _T_49 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_50 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 364:31]
  wire  _T_54 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_147 = _T_54 ? 64'h0 : _GEN_27; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_188 = _T_49 ? _GEN_27 : _GEN_147; // @[Conditional.scala 39:67]
  wire  _GEN_221 = _T_38 & _T_40; // @[PhiNode.scala 341:23]
  wire  _GEN_222 = _GEN_221 & enable_R_control; // @[PhiNode.scala 341:23]
  wire  _GEN_223 = _GEN_222 & _T_42; // @[PhiNode.scala 341:23]
  wire  _GEN_227 = ~enable_R_control; // @[PhiNode.scala 357:19]
  wire  _GEN_228 = _GEN_221 & _GEN_227; // @[PhiNode.scala 357:19]
  assign io_enable_ready = ~enable_valid_R; // @[PhiNode.scala 245:19]
  assign io_InData_0_ready = ~in_data_valid_R_0; // @[PhiNode.scala 253:24]
  assign io_InData_1_ready = ~in_data_valid_R_1; // @[PhiNode.scala 253:24]
  assign io_Mask_ready = ~mask_valid_R; // @[PhiNode.scala 238:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 322:21]
  assign io_Out_0_bits_data = _T_38 ? _GEN_27 : _GEN_188; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 322:21]
  assign io_Out_1_bits_data = _T_38 ? _GEN_27 : _GEN_188; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[4:0];
  _RAND_3 = {2{`RANDOM}};
  in_data_R_1_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_R_control = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enable_valid_R = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mask_R = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  mask_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fire_R_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  guard_index = _RAND_15[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_14) begin
      in_data_R_0_taskID <= io_InData_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else if (_T_38) begin
      if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_R_1_taskID <= 5'h0;
      end else if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_R_1_taskID <= 5'h0;
      end else if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_16) begin
      in_data_R_1_taskID <= io_InData_1_bits_taskID;
    end
    if (reset) begin
      in_data_R_1_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_16) begin
      in_data_R_1_data <= io_InData_1_bits_data;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      in_data_valid_R_0 <= _GEN_11;
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_11;
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else if (_T_38) begin
      in_data_valid_R_1 <= _GEN_15;
    end else if (_T_49) begin
      if (_T_50) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else begin
      in_data_valid_R_1 <= _GEN_15;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_38) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_38) begin
      enable_valid_R <= _GEN_7;
    end else if (_T_49) begin
      if (_T_50) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else begin
      enable_valid_R <= _GEN_7;
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else if (_T_38) begin
      if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_49) begin
      if (_T_50) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_10) begin
      mask_R <= io_Mask_bits;
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else if (_T_38) begin
      mask_valid_R <= _GEN_3;
    end else if (_T_49) begin
      if (_T_50) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else begin
      mask_valid_R <= _GEN_3;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_38) begin
      if (_T_40) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_49) begin
      if (_T_50) begin
        state <= 2'h0;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      out_valid_R_0 <= _GEN_107;
    end else if (_T_17) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_38) begin
      out_valid_R_1 <= _GEN_108;
    end else if (_T_18) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else if (_T_38) begin
      fire_R_0 <= _GEN_16;
    end else if (_T_49) begin
      if (_T_50) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else begin
      fire_R_0 <= _GEN_16;
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else if (_T_38) begin
      fire_R_1 <= _GEN_18;
    end else if (_T_49) begin
      if (_T_50) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else if (_T_54) begin
      if (_T_50) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else begin
      fire_R_1 <= _GEN_18;
    end
    if (reset) begin
      guard_index <= 6'h0;
    end else if (_T_33) begin
      guard_index <= _T_37;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_223 & _T_44) begin
          $fwrite(32'h80000002,"[DEBUG] [Bbgemm] [TID->%d] [PHI] phiindvars_iv823 Produced value: %d, correct value: %d\n",_GEN_26,_GEN_27,_GEN_91); // @[PhiNode.scala 341:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_222 & _T_44) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv823] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_102,enable_R_control,_GEN_27,cycleCount); // @[PhiNode.scala 350:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_228 & _T_44) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv823] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_102,enable_R_control,_GEN_27,cycleCount); // @[PhiNode.scala 357:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_2(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  state; // @[BranchNode.scala 588:22]
  wire  _T_11 = ~state; // @[Conditional.scala 37:30]
  wire  _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_16 = ~reset; // @[BranchNode.scala 616:17]
  wire  _GEN_8 = enable_valid_R | state; // @[BranchNode.scala 611:46]
  wire  _GEN_10 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 611:46]
  wire  _T_18 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_19 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_20 = _T_18 | _T_19; // @[HandShaking.scala 725:29]
  wire  _GEN_31 = _T_11 & enable_valid_R; // @[BranchNode.scala 616:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = _T_11 ? _GEN_10 : out_valid_R_0; // @[HandShaking.scala 630:21 BranchNode.scala 614:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 607:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 607:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_control <= 1'h0;
      end else if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_20) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (enable_valid_R) begin
        out_valid_R_0 <= _T_14;
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_11) begin
      state <= _GEN_8;
    end else if (state) begin
      if (_T_20) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [UBR] [br_4] [Out: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,cycleCount); // @[BranchNode.scala 616:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [63:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] in_data_R_0_taskID; // @[PhiNode.scala 203:26]
  reg [4:0] in_data_R_1_taskID; // @[PhiNode.scala 203:26]
  reg [63:0] in_data_R_1_data; // @[PhiNode.scala 203:26]
  reg  in_data_valid_R_0; // @[PhiNode.scala 204:32]
  reg  in_data_valid_R_1; // @[PhiNode.scala 204:32]
  reg  enable_R_control; // @[PhiNode.scala 207:25]
  reg  enable_valid_R; // @[PhiNode.scala 208:31]
  reg [1:0] mask_R; // @[PhiNode.scala 211:23]
  reg  mask_valid_R; // @[PhiNode.scala 212:29]
  reg [1:0] state; // @[PhiNode.scala 216:22]
  reg  out_valid_R_0; // @[PhiNode.scala 219:49]
  reg  out_valid_R_1; // @[PhiNode.scala 219:49]
  reg  fire_R_0; // @[PhiNode.scala 221:44]
  reg  fire_R_1; // @[PhiNode.scala 221:44]
  wire  _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_10 | mask_valid_R; // @[PhiNode.scala 239:24]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_12 | enable_valid_R; // @[PhiNode.scala 246:26]
  wire  _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 254:29]
  wire  _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 254:29]
  wire [1:0] _T_19 = {mask_R[0],mask_R[1]}; // @[Cat.scala 29:58]
  wire  sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  wire  _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_16 = _T_20 | fire_R_0; // @[PhiNode.scala 276:26]
  wire  _GEN_17 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 276:26]
  wire  _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = _T_21 | fire_R_1; // @[PhiNode.scala 276:26]
  wire  _GEN_19 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 276:26]
  wire  fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 283:74]
  wire  fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 283:74]
  wire [63:0] _GEN_27 = sel ? in_data_R_1_data : 64'h0; // @[PhiNode.scala 312:12]
  wire  _T_41 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_42 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 286:30]
  wire  _T_43 = enable_valid_R & _T_42; // @[PhiNode.scala 327:27]
  reg [9:0] guard_index; // @[Counter.scala 29:33]
  wire [63:0] _GEN_29 = 10'h1 == guard_index ? 64'h1 : 64'h0; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_30 = 10'h2 == guard_index ? 64'h2 : _GEN_29; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_31 = 10'h3 == guard_index ? 64'h3 : _GEN_30; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_32 = 10'h4 == guard_index ? 64'h4 : _GEN_31; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_33 = 10'h5 == guard_index ? 64'h5 : _GEN_32; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_34 = 10'h6 == guard_index ? 64'h6 : _GEN_33; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_35 = 10'h7 == guard_index ? 64'h7 : _GEN_34; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_36 = 10'h8 == guard_index ? 64'h8 : _GEN_35; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_37 = 10'h9 == guard_index ? 64'h9 : _GEN_36; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_38 = 10'ha == guard_index ? 64'ha : _GEN_37; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_39 = 10'hb == guard_index ? 64'hb : _GEN_38; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_40 = 10'hc == guard_index ? 64'hc : _GEN_39; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_41 = 10'hd == guard_index ? 64'hd : _GEN_40; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_42 = 10'he == guard_index ? 64'he : _GEN_41; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_43 = 10'hf == guard_index ? 64'hf : _GEN_42; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_44 = 10'h10 == guard_index ? 64'h0 : _GEN_43; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_45 = 10'h11 == guard_index ? 64'h1 : _GEN_44; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_46 = 10'h12 == guard_index ? 64'h2 : _GEN_45; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_47 = 10'h13 == guard_index ? 64'h3 : _GEN_46; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_48 = 10'h14 == guard_index ? 64'h4 : _GEN_47; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_49 = 10'h15 == guard_index ? 64'h5 : _GEN_48; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_50 = 10'h16 == guard_index ? 64'h6 : _GEN_49; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_51 = 10'h17 == guard_index ? 64'h7 : _GEN_50; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_52 = 10'h18 == guard_index ? 64'h8 : _GEN_51; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_53 = 10'h19 == guard_index ? 64'h9 : _GEN_52; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_54 = 10'h1a == guard_index ? 64'ha : _GEN_53; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_55 = 10'h1b == guard_index ? 64'hb : _GEN_54; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_56 = 10'h1c == guard_index ? 64'hc : _GEN_55; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_57 = 10'h1d == guard_index ? 64'hd : _GEN_56; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_58 = 10'h1e == guard_index ? 64'he : _GEN_57; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_59 = 10'h1f == guard_index ? 64'hf : _GEN_58; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_60 = 10'h20 == guard_index ? 64'h0 : _GEN_59; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_61 = 10'h21 == guard_index ? 64'h1 : _GEN_60; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_62 = 10'h22 == guard_index ? 64'h2 : _GEN_61; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_63 = 10'h23 == guard_index ? 64'h3 : _GEN_62; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_64 = 10'h24 == guard_index ? 64'h4 : _GEN_63; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_65 = 10'h25 == guard_index ? 64'h5 : _GEN_64; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_66 = 10'h26 == guard_index ? 64'h6 : _GEN_65; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_67 = 10'h27 == guard_index ? 64'h7 : _GEN_66; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_68 = 10'h28 == guard_index ? 64'h8 : _GEN_67; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_69 = 10'h29 == guard_index ? 64'h9 : _GEN_68; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_70 = 10'h2a == guard_index ? 64'ha : _GEN_69; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_71 = 10'h2b == guard_index ? 64'hb : _GEN_70; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_72 = 10'h2c == guard_index ? 64'hc : _GEN_71; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_73 = 10'h2d == guard_index ? 64'hd : _GEN_72; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_74 = 10'h2e == guard_index ? 64'he : _GEN_73; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_75 = 10'h2f == guard_index ? 64'hf : _GEN_74; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_76 = 10'h30 == guard_index ? 64'h0 : _GEN_75; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_77 = 10'h31 == guard_index ? 64'h1 : _GEN_76; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_78 = 10'h32 == guard_index ? 64'h2 : _GEN_77; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_79 = 10'h33 == guard_index ? 64'h3 : _GEN_78; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_80 = 10'h34 == guard_index ? 64'h4 : _GEN_79; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_81 = 10'h35 == guard_index ? 64'h5 : _GEN_80; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_82 = 10'h36 == guard_index ? 64'h6 : _GEN_81; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_83 = 10'h37 == guard_index ? 64'h7 : _GEN_82; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_84 = 10'h38 == guard_index ? 64'h8 : _GEN_83; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_85 = 10'h39 == guard_index ? 64'h9 : _GEN_84; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_86 = 10'h3a == guard_index ? 64'ha : _GEN_85; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_87 = 10'h3b == guard_index ? 64'hb : _GEN_86; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_88 = 10'h3c == guard_index ? 64'hc : _GEN_87; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_89 = 10'h3d == guard_index ? 64'hd : _GEN_88; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_90 = 10'h3e == guard_index ? 64'he : _GEN_89; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_91 = 10'h3f == guard_index ? 64'hf : _GEN_90; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_92 = 10'h40 == guard_index ? 64'h0 : _GEN_91; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_93 = 10'h41 == guard_index ? 64'h1 : _GEN_92; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_94 = 10'h42 == guard_index ? 64'h2 : _GEN_93; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_95 = 10'h43 == guard_index ? 64'h3 : _GEN_94; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_96 = 10'h44 == guard_index ? 64'h4 : _GEN_95; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_97 = 10'h45 == guard_index ? 64'h5 : _GEN_96; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_98 = 10'h46 == guard_index ? 64'h6 : _GEN_97; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_99 = 10'h47 == guard_index ? 64'h7 : _GEN_98; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_100 = 10'h48 == guard_index ? 64'h8 : _GEN_99; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_101 = 10'h49 == guard_index ? 64'h9 : _GEN_100; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_102 = 10'h4a == guard_index ? 64'ha : _GEN_101; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_103 = 10'h4b == guard_index ? 64'hb : _GEN_102; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_104 = 10'h4c == guard_index ? 64'hc : _GEN_103; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_105 = 10'h4d == guard_index ? 64'hd : _GEN_104; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_106 = 10'h4e == guard_index ? 64'he : _GEN_105; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_107 = 10'h4f == guard_index ? 64'hf : _GEN_106; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_108 = 10'h50 == guard_index ? 64'h0 : _GEN_107; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_109 = 10'h51 == guard_index ? 64'h1 : _GEN_108; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_110 = 10'h52 == guard_index ? 64'h2 : _GEN_109; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_111 = 10'h53 == guard_index ? 64'h3 : _GEN_110; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_112 = 10'h54 == guard_index ? 64'h4 : _GEN_111; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_113 = 10'h55 == guard_index ? 64'h5 : _GEN_112; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_114 = 10'h56 == guard_index ? 64'h6 : _GEN_113; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_115 = 10'h57 == guard_index ? 64'h7 : _GEN_114; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_116 = 10'h58 == guard_index ? 64'h8 : _GEN_115; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_117 = 10'h59 == guard_index ? 64'h9 : _GEN_116; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_118 = 10'h5a == guard_index ? 64'ha : _GEN_117; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_119 = 10'h5b == guard_index ? 64'hb : _GEN_118; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_120 = 10'h5c == guard_index ? 64'hc : _GEN_119; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_121 = 10'h5d == guard_index ? 64'hd : _GEN_120; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_122 = 10'h5e == guard_index ? 64'he : _GEN_121; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_123 = 10'h5f == guard_index ? 64'hf : _GEN_122; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_124 = 10'h60 == guard_index ? 64'h0 : _GEN_123; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_125 = 10'h61 == guard_index ? 64'h1 : _GEN_124; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_126 = 10'h62 == guard_index ? 64'h2 : _GEN_125; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_127 = 10'h63 == guard_index ? 64'h3 : _GEN_126; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_128 = 10'h64 == guard_index ? 64'h4 : _GEN_127; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_129 = 10'h65 == guard_index ? 64'h5 : _GEN_128; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_130 = 10'h66 == guard_index ? 64'h6 : _GEN_129; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_131 = 10'h67 == guard_index ? 64'h7 : _GEN_130; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_132 = 10'h68 == guard_index ? 64'h8 : _GEN_131; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_133 = 10'h69 == guard_index ? 64'h9 : _GEN_132; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_134 = 10'h6a == guard_index ? 64'ha : _GEN_133; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_135 = 10'h6b == guard_index ? 64'hb : _GEN_134; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_136 = 10'h6c == guard_index ? 64'hc : _GEN_135; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_137 = 10'h6d == guard_index ? 64'hd : _GEN_136; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_138 = 10'h6e == guard_index ? 64'he : _GEN_137; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_139 = 10'h6f == guard_index ? 64'hf : _GEN_138; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_140 = 10'h70 == guard_index ? 64'h0 : _GEN_139; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_141 = 10'h71 == guard_index ? 64'h1 : _GEN_140; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_142 = 10'h72 == guard_index ? 64'h2 : _GEN_141; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_143 = 10'h73 == guard_index ? 64'h3 : _GEN_142; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_144 = 10'h74 == guard_index ? 64'h4 : _GEN_143; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_145 = 10'h75 == guard_index ? 64'h5 : _GEN_144; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_146 = 10'h76 == guard_index ? 64'h6 : _GEN_145; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_147 = 10'h77 == guard_index ? 64'h7 : _GEN_146; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_148 = 10'h78 == guard_index ? 64'h8 : _GEN_147; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_149 = 10'h79 == guard_index ? 64'h9 : _GEN_148; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_150 = 10'h7a == guard_index ? 64'ha : _GEN_149; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_151 = 10'h7b == guard_index ? 64'hb : _GEN_150; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_152 = 10'h7c == guard_index ? 64'hc : _GEN_151; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_153 = 10'h7d == guard_index ? 64'hd : _GEN_152; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_154 = 10'h7e == guard_index ? 64'he : _GEN_153; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_155 = 10'h7f == guard_index ? 64'hf : _GEN_154; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_156 = 10'h80 == guard_index ? 64'h0 : _GEN_155; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_157 = 10'h81 == guard_index ? 64'h1 : _GEN_156; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_158 = 10'h82 == guard_index ? 64'h2 : _GEN_157; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_159 = 10'h83 == guard_index ? 64'h3 : _GEN_158; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_160 = 10'h84 == guard_index ? 64'h4 : _GEN_159; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_161 = 10'h85 == guard_index ? 64'h5 : _GEN_160; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_162 = 10'h86 == guard_index ? 64'h6 : _GEN_161; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_163 = 10'h87 == guard_index ? 64'h7 : _GEN_162; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_164 = 10'h88 == guard_index ? 64'h8 : _GEN_163; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_165 = 10'h89 == guard_index ? 64'h9 : _GEN_164; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_166 = 10'h8a == guard_index ? 64'ha : _GEN_165; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_167 = 10'h8b == guard_index ? 64'hb : _GEN_166; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_168 = 10'h8c == guard_index ? 64'hc : _GEN_167; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_169 = 10'h8d == guard_index ? 64'hd : _GEN_168; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_170 = 10'h8e == guard_index ? 64'he : _GEN_169; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_171 = 10'h8f == guard_index ? 64'hf : _GEN_170; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_172 = 10'h90 == guard_index ? 64'h0 : _GEN_171; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_173 = 10'h91 == guard_index ? 64'h1 : _GEN_172; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_174 = 10'h92 == guard_index ? 64'h2 : _GEN_173; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_175 = 10'h93 == guard_index ? 64'h3 : _GEN_174; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_176 = 10'h94 == guard_index ? 64'h4 : _GEN_175; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_177 = 10'h95 == guard_index ? 64'h5 : _GEN_176; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_178 = 10'h96 == guard_index ? 64'h6 : _GEN_177; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_179 = 10'h97 == guard_index ? 64'h7 : _GEN_178; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_180 = 10'h98 == guard_index ? 64'h8 : _GEN_179; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_181 = 10'h99 == guard_index ? 64'h9 : _GEN_180; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_182 = 10'h9a == guard_index ? 64'ha : _GEN_181; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_183 = 10'h9b == guard_index ? 64'hb : _GEN_182; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_184 = 10'h9c == guard_index ? 64'hc : _GEN_183; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_185 = 10'h9d == guard_index ? 64'hd : _GEN_184; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_186 = 10'h9e == guard_index ? 64'he : _GEN_185; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_187 = 10'h9f == guard_index ? 64'hf : _GEN_186; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_188 = 10'ha0 == guard_index ? 64'h0 : _GEN_187; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_189 = 10'ha1 == guard_index ? 64'h1 : _GEN_188; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_190 = 10'ha2 == guard_index ? 64'h2 : _GEN_189; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_191 = 10'ha3 == guard_index ? 64'h3 : _GEN_190; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_192 = 10'ha4 == guard_index ? 64'h4 : _GEN_191; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_193 = 10'ha5 == guard_index ? 64'h5 : _GEN_192; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_194 = 10'ha6 == guard_index ? 64'h6 : _GEN_193; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_195 = 10'ha7 == guard_index ? 64'h7 : _GEN_194; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_196 = 10'ha8 == guard_index ? 64'h8 : _GEN_195; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_197 = 10'ha9 == guard_index ? 64'h9 : _GEN_196; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_198 = 10'haa == guard_index ? 64'ha : _GEN_197; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_199 = 10'hab == guard_index ? 64'hb : _GEN_198; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_200 = 10'hac == guard_index ? 64'hc : _GEN_199; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_201 = 10'had == guard_index ? 64'hd : _GEN_200; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_202 = 10'hae == guard_index ? 64'he : _GEN_201; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_203 = 10'haf == guard_index ? 64'hf : _GEN_202; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_204 = 10'hb0 == guard_index ? 64'h0 : _GEN_203; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_205 = 10'hb1 == guard_index ? 64'h1 : _GEN_204; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_206 = 10'hb2 == guard_index ? 64'h2 : _GEN_205; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_207 = 10'hb3 == guard_index ? 64'h3 : _GEN_206; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_208 = 10'hb4 == guard_index ? 64'h4 : _GEN_207; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_209 = 10'hb5 == guard_index ? 64'h5 : _GEN_208; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_210 = 10'hb6 == guard_index ? 64'h6 : _GEN_209; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_211 = 10'hb7 == guard_index ? 64'h7 : _GEN_210; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_212 = 10'hb8 == guard_index ? 64'h8 : _GEN_211; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_213 = 10'hb9 == guard_index ? 64'h9 : _GEN_212; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_214 = 10'hba == guard_index ? 64'ha : _GEN_213; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_215 = 10'hbb == guard_index ? 64'hb : _GEN_214; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_216 = 10'hbc == guard_index ? 64'hc : _GEN_215; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_217 = 10'hbd == guard_index ? 64'hd : _GEN_216; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_218 = 10'hbe == guard_index ? 64'he : _GEN_217; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_219 = 10'hbf == guard_index ? 64'hf : _GEN_218; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_220 = 10'hc0 == guard_index ? 64'h0 : _GEN_219; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_221 = 10'hc1 == guard_index ? 64'h1 : _GEN_220; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_222 = 10'hc2 == guard_index ? 64'h2 : _GEN_221; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_223 = 10'hc3 == guard_index ? 64'h3 : _GEN_222; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_224 = 10'hc4 == guard_index ? 64'h4 : _GEN_223; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_225 = 10'hc5 == guard_index ? 64'h5 : _GEN_224; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_226 = 10'hc6 == guard_index ? 64'h6 : _GEN_225; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_227 = 10'hc7 == guard_index ? 64'h7 : _GEN_226; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_228 = 10'hc8 == guard_index ? 64'h8 : _GEN_227; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_229 = 10'hc9 == guard_index ? 64'h9 : _GEN_228; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_230 = 10'hca == guard_index ? 64'ha : _GEN_229; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_231 = 10'hcb == guard_index ? 64'hb : _GEN_230; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_232 = 10'hcc == guard_index ? 64'hc : _GEN_231; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_233 = 10'hcd == guard_index ? 64'hd : _GEN_232; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_234 = 10'hce == guard_index ? 64'he : _GEN_233; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_235 = 10'hcf == guard_index ? 64'hf : _GEN_234; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_236 = 10'hd0 == guard_index ? 64'h0 : _GEN_235; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_237 = 10'hd1 == guard_index ? 64'h1 : _GEN_236; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_238 = 10'hd2 == guard_index ? 64'h2 : _GEN_237; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_239 = 10'hd3 == guard_index ? 64'h3 : _GEN_238; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_240 = 10'hd4 == guard_index ? 64'h4 : _GEN_239; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_241 = 10'hd5 == guard_index ? 64'h5 : _GEN_240; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_242 = 10'hd6 == guard_index ? 64'h6 : _GEN_241; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_243 = 10'hd7 == guard_index ? 64'h7 : _GEN_242; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_244 = 10'hd8 == guard_index ? 64'h8 : _GEN_243; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_245 = 10'hd9 == guard_index ? 64'h9 : _GEN_244; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_246 = 10'hda == guard_index ? 64'ha : _GEN_245; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_247 = 10'hdb == guard_index ? 64'hb : _GEN_246; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_248 = 10'hdc == guard_index ? 64'hc : _GEN_247; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_249 = 10'hdd == guard_index ? 64'hd : _GEN_248; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_250 = 10'hde == guard_index ? 64'he : _GEN_249; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_251 = 10'hdf == guard_index ? 64'hf : _GEN_250; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_252 = 10'he0 == guard_index ? 64'h0 : _GEN_251; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_253 = 10'he1 == guard_index ? 64'h1 : _GEN_252; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_254 = 10'he2 == guard_index ? 64'h2 : _GEN_253; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_255 = 10'he3 == guard_index ? 64'h3 : _GEN_254; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_256 = 10'he4 == guard_index ? 64'h4 : _GEN_255; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_257 = 10'he5 == guard_index ? 64'h5 : _GEN_256; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_258 = 10'he6 == guard_index ? 64'h6 : _GEN_257; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_259 = 10'he7 == guard_index ? 64'h7 : _GEN_258; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_260 = 10'he8 == guard_index ? 64'h8 : _GEN_259; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_261 = 10'he9 == guard_index ? 64'h9 : _GEN_260; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_262 = 10'hea == guard_index ? 64'ha : _GEN_261; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_263 = 10'heb == guard_index ? 64'hb : _GEN_262; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_264 = 10'hec == guard_index ? 64'hc : _GEN_263; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_265 = 10'hed == guard_index ? 64'hd : _GEN_264; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_266 = 10'hee == guard_index ? 64'he : _GEN_265; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_267 = 10'hef == guard_index ? 64'hf : _GEN_266; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_268 = 10'hf0 == guard_index ? 64'h0 : _GEN_267; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_269 = 10'hf1 == guard_index ? 64'h1 : _GEN_268; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_270 = 10'hf2 == guard_index ? 64'h2 : _GEN_269; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_271 = 10'hf3 == guard_index ? 64'h3 : _GEN_270; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_272 = 10'hf4 == guard_index ? 64'h4 : _GEN_271; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_273 = 10'hf5 == guard_index ? 64'h5 : _GEN_272; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_274 = 10'hf6 == guard_index ? 64'h6 : _GEN_273; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_275 = 10'hf7 == guard_index ? 64'h7 : _GEN_274; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_276 = 10'hf8 == guard_index ? 64'h8 : _GEN_275; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_277 = 10'hf9 == guard_index ? 64'h9 : _GEN_276; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_278 = 10'hfa == guard_index ? 64'ha : _GEN_277; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_279 = 10'hfb == guard_index ? 64'hb : _GEN_278; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_280 = 10'hfc == guard_index ? 64'hc : _GEN_279; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_281 = 10'hfd == guard_index ? 64'hd : _GEN_280; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_282 = 10'hfe == guard_index ? 64'he : _GEN_281; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_283 = 10'hff == guard_index ? 64'hf : _GEN_282; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_284 = 10'h100 == guard_index ? 64'h0 : _GEN_283; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_285 = 10'h101 == guard_index ? 64'h1 : _GEN_284; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_286 = 10'h102 == guard_index ? 64'h2 : _GEN_285; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_287 = 10'h103 == guard_index ? 64'h3 : _GEN_286; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_288 = 10'h104 == guard_index ? 64'h4 : _GEN_287; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_289 = 10'h105 == guard_index ? 64'h5 : _GEN_288; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_290 = 10'h106 == guard_index ? 64'h6 : _GEN_289; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_291 = 10'h107 == guard_index ? 64'h7 : _GEN_290; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_292 = 10'h108 == guard_index ? 64'h8 : _GEN_291; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_293 = 10'h109 == guard_index ? 64'h9 : _GEN_292; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_294 = 10'h10a == guard_index ? 64'ha : _GEN_293; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_295 = 10'h10b == guard_index ? 64'hb : _GEN_294; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_296 = 10'h10c == guard_index ? 64'hc : _GEN_295; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_297 = 10'h10d == guard_index ? 64'hd : _GEN_296; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_298 = 10'h10e == guard_index ? 64'he : _GEN_297; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_299 = 10'h10f == guard_index ? 64'hf : _GEN_298; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_300 = 10'h110 == guard_index ? 64'h0 : _GEN_299; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_301 = 10'h111 == guard_index ? 64'h1 : _GEN_300; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_302 = 10'h112 == guard_index ? 64'h2 : _GEN_301; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_303 = 10'h113 == guard_index ? 64'h3 : _GEN_302; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_304 = 10'h114 == guard_index ? 64'h4 : _GEN_303; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_305 = 10'h115 == guard_index ? 64'h5 : _GEN_304; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_306 = 10'h116 == guard_index ? 64'h6 : _GEN_305; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_307 = 10'h117 == guard_index ? 64'h7 : _GEN_306; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_308 = 10'h118 == guard_index ? 64'h8 : _GEN_307; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_309 = 10'h119 == guard_index ? 64'h9 : _GEN_308; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_310 = 10'h11a == guard_index ? 64'ha : _GEN_309; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_311 = 10'h11b == guard_index ? 64'hb : _GEN_310; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_312 = 10'h11c == guard_index ? 64'hc : _GEN_311; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_313 = 10'h11d == guard_index ? 64'hd : _GEN_312; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_314 = 10'h11e == guard_index ? 64'he : _GEN_313; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_315 = 10'h11f == guard_index ? 64'hf : _GEN_314; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_316 = 10'h120 == guard_index ? 64'h0 : _GEN_315; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_317 = 10'h121 == guard_index ? 64'h1 : _GEN_316; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_318 = 10'h122 == guard_index ? 64'h2 : _GEN_317; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_319 = 10'h123 == guard_index ? 64'h3 : _GEN_318; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_320 = 10'h124 == guard_index ? 64'h4 : _GEN_319; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_321 = 10'h125 == guard_index ? 64'h5 : _GEN_320; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_322 = 10'h126 == guard_index ? 64'h6 : _GEN_321; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_323 = 10'h127 == guard_index ? 64'h7 : _GEN_322; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_324 = 10'h128 == guard_index ? 64'h8 : _GEN_323; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_325 = 10'h129 == guard_index ? 64'h9 : _GEN_324; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_326 = 10'h12a == guard_index ? 64'ha : _GEN_325; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_327 = 10'h12b == guard_index ? 64'hb : _GEN_326; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_328 = 10'h12c == guard_index ? 64'hc : _GEN_327; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_329 = 10'h12d == guard_index ? 64'hd : _GEN_328; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_330 = 10'h12e == guard_index ? 64'he : _GEN_329; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_331 = 10'h12f == guard_index ? 64'hf : _GEN_330; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_332 = 10'h130 == guard_index ? 64'h0 : _GEN_331; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_333 = 10'h131 == guard_index ? 64'h1 : _GEN_332; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_334 = 10'h132 == guard_index ? 64'h2 : _GEN_333; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_335 = 10'h133 == guard_index ? 64'h3 : _GEN_334; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_336 = 10'h134 == guard_index ? 64'h4 : _GEN_335; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_337 = 10'h135 == guard_index ? 64'h5 : _GEN_336; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_338 = 10'h136 == guard_index ? 64'h6 : _GEN_337; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_339 = 10'h137 == guard_index ? 64'h7 : _GEN_338; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_340 = 10'h138 == guard_index ? 64'h8 : _GEN_339; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_341 = 10'h139 == guard_index ? 64'h9 : _GEN_340; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_342 = 10'h13a == guard_index ? 64'ha : _GEN_341; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_343 = 10'h13b == guard_index ? 64'hb : _GEN_342; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_344 = 10'h13c == guard_index ? 64'hc : _GEN_343; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_345 = 10'h13d == guard_index ? 64'hd : _GEN_344; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_346 = 10'h13e == guard_index ? 64'he : _GEN_345; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_347 = 10'h13f == guard_index ? 64'hf : _GEN_346; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_348 = 10'h140 == guard_index ? 64'h0 : _GEN_347; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_349 = 10'h141 == guard_index ? 64'h1 : _GEN_348; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_350 = 10'h142 == guard_index ? 64'h2 : _GEN_349; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_351 = 10'h143 == guard_index ? 64'h3 : _GEN_350; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_352 = 10'h144 == guard_index ? 64'h4 : _GEN_351; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_353 = 10'h145 == guard_index ? 64'h5 : _GEN_352; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_354 = 10'h146 == guard_index ? 64'h6 : _GEN_353; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_355 = 10'h147 == guard_index ? 64'h7 : _GEN_354; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_356 = 10'h148 == guard_index ? 64'h8 : _GEN_355; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_357 = 10'h149 == guard_index ? 64'h9 : _GEN_356; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_358 = 10'h14a == guard_index ? 64'ha : _GEN_357; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_359 = 10'h14b == guard_index ? 64'hb : _GEN_358; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_360 = 10'h14c == guard_index ? 64'hc : _GEN_359; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_361 = 10'h14d == guard_index ? 64'hd : _GEN_360; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_362 = 10'h14e == guard_index ? 64'he : _GEN_361; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_363 = 10'h14f == guard_index ? 64'hf : _GEN_362; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_364 = 10'h150 == guard_index ? 64'h0 : _GEN_363; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_365 = 10'h151 == guard_index ? 64'h1 : _GEN_364; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_366 = 10'h152 == guard_index ? 64'h2 : _GEN_365; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_367 = 10'h153 == guard_index ? 64'h3 : _GEN_366; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_368 = 10'h154 == guard_index ? 64'h4 : _GEN_367; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_369 = 10'h155 == guard_index ? 64'h5 : _GEN_368; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_370 = 10'h156 == guard_index ? 64'h6 : _GEN_369; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_371 = 10'h157 == guard_index ? 64'h7 : _GEN_370; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_372 = 10'h158 == guard_index ? 64'h8 : _GEN_371; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_373 = 10'h159 == guard_index ? 64'h9 : _GEN_372; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_374 = 10'h15a == guard_index ? 64'ha : _GEN_373; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_375 = 10'h15b == guard_index ? 64'hb : _GEN_374; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_376 = 10'h15c == guard_index ? 64'hc : _GEN_375; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_377 = 10'h15d == guard_index ? 64'hd : _GEN_376; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_378 = 10'h15e == guard_index ? 64'he : _GEN_377; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_379 = 10'h15f == guard_index ? 64'hf : _GEN_378; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_380 = 10'h160 == guard_index ? 64'h0 : _GEN_379; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_381 = 10'h161 == guard_index ? 64'h1 : _GEN_380; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_382 = 10'h162 == guard_index ? 64'h2 : _GEN_381; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_383 = 10'h163 == guard_index ? 64'h3 : _GEN_382; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_384 = 10'h164 == guard_index ? 64'h4 : _GEN_383; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_385 = 10'h165 == guard_index ? 64'h5 : _GEN_384; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_386 = 10'h166 == guard_index ? 64'h6 : _GEN_385; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_387 = 10'h167 == guard_index ? 64'h7 : _GEN_386; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_388 = 10'h168 == guard_index ? 64'h8 : _GEN_387; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_389 = 10'h169 == guard_index ? 64'h9 : _GEN_388; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_390 = 10'h16a == guard_index ? 64'ha : _GEN_389; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_391 = 10'h16b == guard_index ? 64'hb : _GEN_390; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_392 = 10'h16c == guard_index ? 64'hc : _GEN_391; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_393 = 10'h16d == guard_index ? 64'hd : _GEN_392; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_394 = 10'h16e == guard_index ? 64'he : _GEN_393; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_395 = 10'h16f == guard_index ? 64'hf : _GEN_394; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_396 = 10'h170 == guard_index ? 64'h0 : _GEN_395; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_397 = 10'h171 == guard_index ? 64'h1 : _GEN_396; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_398 = 10'h172 == guard_index ? 64'h2 : _GEN_397; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_399 = 10'h173 == guard_index ? 64'h3 : _GEN_398; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_400 = 10'h174 == guard_index ? 64'h4 : _GEN_399; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_401 = 10'h175 == guard_index ? 64'h5 : _GEN_400; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_402 = 10'h176 == guard_index ? 64'h6 : _GEN_401; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_403 = 10'h177 == guard_index ? 64'h7 : _GEN_402; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_404 = 10'h178 == guard_index ? 64'h8 : _GEN_403; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_405 = 10'h179 == guard_index ? 64'h9 : _GEN_404; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_406 = 10'h17a == guard_index ? 64'ha : _GEN_405; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_407 = 10'h17b == guard_index ? 64'hb : _GEN_406; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_408 = 10'h17c == guard_index ? 64'hc : _GEN_407; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_409 = 10'h17d == guard_index ? 64'hd : _GEN_408; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_410 = 10'h17e == guard_index ? 64'he : _GEN_409; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_411 = 10'h17f == guard_index ? 64'hf : _GEN_410; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_412 = 10'h180 == guard_index ? 64'h0 : _GEN_411; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_413 = 10'h181 == guard_index ? 64'h1 : _GEN_412; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_414 = 10'h182 == guard_index ? 64'h2 : _GEN_413; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_415 = 10'h183 == guard_index ? 64'h3 : _GEN_414; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_416 = 10'h184 == guard_index ? 64'h4 : _GEN_415; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_417 = 10'h185 == guard_index ? 64'h5 : _GEN_416; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_418 = 10'h186 == guard_index ? 64'h6 : _GEN_417; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_419 = 10'h187 == guard_index ? 64'h7 : _GEN_418; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_420 = 10'h188 == guard_index ? 64'h8 : _GEN_419; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_421 = 10'h189 == guard_index ? 64'h9 : _GEN_420; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_422 = 10'h18a == guard_index ? 64'ha : _GEN_421; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_423 = 10'h18b == guard_index ? 64'hb : _GEN_422; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_424 = 10'h18c == guard_index ? 64'hc : _GEN_423; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_425 = 10'h18d == guard_index ? 64'hd : _GEN_424; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_426 = 10'h18e == guard_index ? 64'he : _GEN_425; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_427 = 10'h18f == guard_index ? 64'hf : _GEN_426; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_428 = 10'h190 == guard_index ? 64'h0 : _GEN_427; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_429 = 10'h191 == guard_index ? 64'h1 : _GEN_428; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_430 = 10'h192 == guard_index ? 64'h2 : _GEN_429; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_431 = 10'h193 == guard_index ? 64'h3 : _GEN_430; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_432 = 10'h194 == guard_index ? 64'h4 : _GEN_431; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_433 = 10'h195 == guard_index ? 64'h5 : _GEN_432; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_434 = 10'h196 == guard_index ? 64'h6 : _GEN_433; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_435 = 10'h197 == guard_index ? 64'h7 : _GEN_434; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_436 = 10'h198 == guard_index ? 64'h8 : _GEN_435; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_437 = 10'h199 == guard_index ? 64'h9 : _GEN_436; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_438 = 10'h19a == guard_index ? 64'ha : _GEN_437; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_439 = 10'h19b == guard_index ? 64'hb : _GEN_438; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_440 = 10'h19c == guard_index ? 64'hc : _GEN_439; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_441 = 10'h19d == guard_index ? 64'hd : _GEN_440; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_442 = 10'h19e == guard_index ? 64'he : _GEN_441; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_443 = 10'h19f == guard_index ? 64'hf : _GEN_442; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_444 = 10'h1a0 == guard_index ? 64'h0 : _GEN_443; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_445 = 10'h1a1 == guard_index ? 64'h1 : _GEN_444; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_446 = 10'h1a2 == guard_index ? 64'h2 : _GEN_445; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_447 = 10'h1a3 == guard_index ? 64'h3 : _GEN_446; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_448 = 10'h1a4 == guard_index ? 64'h4 : _GEN_447; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_449 = 10'h1a5 == guard_index ? 64'h5 : _GEN_448; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_450 = 10'h1a6 == guard_index ? 64'h6 : _GEN_449; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_451 = 10'h1a7 == guard_index ? 64'h7 : _GEN_450; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_452 = 10'h1a8 == guard_index ? 64'h8 : _GEN_451; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_453 = 10'h1a9 == guard_index ? 64'h9 : _GEN_452; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_454 = 10'h1aa == guard_index ? 64'ha : _GEN_453; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_455 = 10'h1ab == guard_index ? 64'hb : _GEN_454; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_456 = 10'h1ac == guard_index ? 64'hc : _GEN_455; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_457 = 10'h1ad == guard_index ? 64'hd : _GEN_456; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_458 = 10'h1ae == guard_index ? 64'he : _GEN_457; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_459 = 10'h1af == guard_index ? 64'hf : _GEN_458; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_460 = 10'h1b0 == guard_index ? 64'h0 : _GEN_459; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_461 = 10'h1b1 == guard_index ? 64'h1 : _GEN_460; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_462 = 10'h1b2 == guard_index ? 64'h2 : _GEN_461; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_463 = 10'h1b3 == guard_index ? 64'h3 : _GEN_462; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_464 = 10'h1b4 == guard_index ? 64'h4 : _GEN_463; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_465 = 10'h1b5 == guard_index ? 64'h5 : _GEN_464; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_466 = 10'h1b6 == guard_index ? 64'h6 : _GEN_465; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_467 = 10'h1b7 == guard_index ? 64'h7 : _GEN_466; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_468 = 10'h1b8 == guard_index ? 64'h8 : _GEN_467; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_469 = 10'h1b9 == guard_index ? 64'h9 : _GEN_468; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_470 = 10'h1ba == guard_index ? 64'ha : _GEN_469; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_471 = 10'h1bb == guard_index ? 64'hb : _GEN_470; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_472 = 10'h1bc == guard_index ? 64'hc : _GEN_471; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_473 = 10'h1bd == guard_index ? 64'hd : _GEN_472; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_474 = 10'h1be == guard_index ? 64'he : _GEN_473; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_475 = 10'h1bf == guard_index ? 64'hf : _GEN_474; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_476 = 10'h1c0 == guard_index ? 64'h0 : _GEN_475; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_477 = 10'h1c1 == guard_index ? 64'h1 : _GEN_476; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_478 = 10'h1c2 == guard_index ? 64'h2 : _GEN_477; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_479 = 10'h1c3 == guard_index ? 64'h3 : _GEN_478; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_480 = 10'h1c4 == guard_index ? 64'h4 : _GEN_479; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_481 = 10'h1c5 == guard_index ? 64'h5 : _GEN_480; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_482 = 10'h1c6 == guard_index ? 64'h6 : _GEN_481; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_483 = 10'h1c7 == guard_index ? 64'h7 : _GEN_482; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_484 = 10'h1c8 == guard_index ? 64'h8 : _GEN_483; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_485 = 10'h1c9 == guard_index ? 64'h9 : _GEN_484; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_486 = 10'h1ca == guard_index ? 64'ha : _GEN_485; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_487 = 10'h1cb == guard_index ? 64'hb : _GEN_486; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_488 = 10'h1cc == guard_index ? 64'hc : _GEN_487; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_489 = 10'h1cd == guard_index ? 64'hd : _GEN_488; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_490 = 10'h1ce == guard_index ? 64'he : _GEN_489; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_491 = 10'h1cf == guard_index ? 64'hf : _GEN_490; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_492 = 10'h1d0 == guard_index ? 64'h0 : _GEN_491; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_493 = 10'h1d1 == guard_index ? 64'h1 : _GEN_492; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_494 = 10'h1d2 == guard_index ? 64'h2 : _GEN_493; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_495 = 10'h1d3 == guard_index ? 64'h3 : _GEN_494; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_496 = 10'h1d4 == guard_index ? 64'h4 : _GEN_495; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_497 = 10'h1d5 == guard_index ? 64'h5 : _GEN_496; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_498 = 10'h1d6 == guard_index ? 64'h6 : _GEN_497; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_499 = 10'h1d7 == guard_index ? 64'h7 : _GEN_498; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_500 = 10'h1d8 == guard_index ? 64'h8 : _GEN_499; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_501 = 10'h1d9 == guard_index ? 64'h9 : _GEN_500; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_502 = 10'h1da == guard_index ? 64'ha : _GEN_501; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_503 = 10'h1db == guard_index ? 64'hb : _GEN_502; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_504 = 10'h1dc == guard_index ? 64'hc : _GEN_503; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_505 = 10'h1dd == guard_index ? 64'hd : _GEN_504; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_506 = 10'h1de == guard_index ? 64'he : _GEN_505; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_507 = 10'h1df == guard_index ? 64'hf : _GEN_506; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_508 = 10'h1e0 == guard_index ? 64'h0 : _GEN_507; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_509 = 10'h1e1 == guard_index ? 64'h1 : _GEN_508; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_510 = 10'h1e2 == guard_index ? 64'h2 : _GEN_509; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_511 = 10'h1e3 == guard_index ? 64'h3 : _GEN_510; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_512 = 10'h1e4 == guard_index ? 64'h4 : _GEN_511; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_513 = 10'h1e5 == guard_index ? 64'h5 : _GEN_512; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_514 = 10'h1e6 == guard_index ? 64'h6 : _GEN_513; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_515 = 10'h1e7 == guard_index ? 64'h7 : _GEN_514; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_516 = 10'h1e8 == guard_index ? 64'h8 : _GEN_515; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_517 = 10'h1e9 == guard_index ? 64'h9 : _GEN_516; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_518 = 10'h1ea == guard_index ? 64'ha : _GEN_517; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_519 = 10'h1eb == guard_index ? 64'hb : _GEN_518; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_520 = 10'h1ec == guard_index ? 64'hc : _GEN_519; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_521 = 10'h1ed == guard_index ? 64'hd : _GEN_520; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_522 = 10'h1ee == guard_index ? 64'he : _GEN_521; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_523 = 10'h1ef == guard_index ? 64'hf : _GEN_522; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_524 = 10'h1f0 == guard_index ? 64'h0 : _GEN_523; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_525 = 10'h1f1 == guard_index ? 64'h1 : _GEN_524; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_526 = 10'h1f2 == guard_index ? 64'h2 : _GEN_525; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_527 = 10'h1f3 == guard_index ? 64'h3 : _GEN_526; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_528 = 10'h1f4 == guard_index ? 64'h4 : _GEN_527; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_529 = 10'h1f5 == guard_index ? 64'h5 : _GEN_528; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_530 = 10'h1f6 == guard_index ? 64'h6 : _GEN_529; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_531 = 10'h1f7 == guard_index ? 64'h7 : _GEN_530; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_532 = 10'h1f8 == guard_index ? 64'h8 : _GEN_531; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_533 = 10'h1f9 == guard_index ? 64'h9 : _GEN_532; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_534 = 10'h1fa == guard_index ? 64'ha : _GEN_533; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_535 = 10'h1fb == guard_index ? 64'hb : _GEN_534; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_536 = 10'h1fc == guard_index ? 64'hc : _GEN_535; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_537 = 10'h1fd == guard_index ? 64'hd : _GEN_536; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_538 = 10'h1fe == guard_index ? 64'he : _GEN_537; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_539 = 10'h1ff == guard_index ? 64'hf : _GEN_538; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_540 = 10'h200 == guard_index ? 64'h0 : _GEN_539; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_541 = 10'h201 == guard_index ? 64'h1 : _GEN_540; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_542 = 10'h202 == guard_index ? 64'h2 : _GEN_541; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_543 = 10'h203 == guard_index ? 64'h3 : _GEN_542; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_544 = 10'h204 == guard_index ? 64'h4 : _GEN_543; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_545 = 10'h205 == guard_index ? 64'h5 : _GEN_544; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_546 = 10'h206 == guard_index ? 64'h6 : _GEN_545; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_547 = 10'h207 == guard_index ? 64'h7 : _GEN_546; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_548 = 10'h208 == guard_index ? 64'h8 : _GEN_547; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_549 = 10'h209 == guard_index ? 64'h9 : _GEN_548; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_550 = 10'h20a == guard_index ? 64'ha : _GEN_549; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_551 = 10'h20b == guard_index ? 64'hb : _GEN_550; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_552 = 10'h20c == guard_index ? 64'hc : _GEN_551; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_553 = 10'h20d == guard_index ? 64'hd : _GEN_552; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_554 = 10'h20e == guard_index ? 64'he : _GEN_553; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_555 = 10'h20f == guard_index ? 64'hf : _GEN_554; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_556 = 10'h210 == guard_index ? 64'h0 : _GEN_555; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_557 = 10'h211 == guard_index ? 64'h1 : _GEN_556; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_558 = 10'h212 == guard_index ? 64'h2 : _GEN_557; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_559 = 10'h213 == guard_index ? 64'h3 : _GEN_558; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_560 = 10'h214 == guard_index ? 64'h4 : _GEN_559; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_561 = 10'h215 == guard_index ? 64'h5 : _GEN_560; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_562 = 10'h216 == guard_index ? 64'h6 : _GEN_561; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_563 = 10'h217 == guard_index ? 64'h7 : _GEN_562; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_564 = 10'h218 == guard_index ? 64'h8 : _GEN_563; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_565 = 10'h219 == guard_index ? 64'h9 : _GEN_564; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_566 = 10'h21a == guard_index ? 64'ha : _GEN_565; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_567 = 10'h21b == guard_index ? 64'hb : _GEN_566; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_568 = 10'h21c == guard_index ? 64'hc : _GEN_567; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_569 = 10'h21d == guard_index ? 64'hd : _GEN_568; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_570 = 10'h21e == guard_index ? 64'he : _GEN_569; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_571 = 10'h21f == guard_index ? 64'hf : _GEN_570; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_572 = 10'h220 == guard_index ? 64'h0 : _GEN_571; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_573 = 10'h221 == guard_index ? 64'h1 : _GEN_572; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_574 = 10'h222 == guard_index ? 64'h2 : _GEN_573; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_575 = 10'h223 == guard_index ? 64'h3 : _GEN_574; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_576 = 10'h224 == guard_index ? 64'h4 : _GEN_575; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_577 = 10'h225 == guard_index ? 64'h5 : _GEN_576; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_578 = 10'h226 == guard_index ? 64'h6 : _GEN_577; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_579 = 10'h227 == guard_index ? 64'h7 : _GEN_578; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_580 = 10'h228 == guard_index ? 64'h8 : _GEN_579; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_581 = 10'h229 == guard_index ? 64'h9 : _GEN_580; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_582 = 10'h22a == guard_index ? 64'ha : _GEN_581; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_583 = 10'h22b == guard_index ? 64'hb : _GEN_582; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_584 = 10'h22c == guard_index ? 64'hc : _GEN_583; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_585 = 10'h22d == guard_index ? 64'hd : _GEN_584; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_586 = 10'h22e == guard_index ? 64'he : _GEN_585; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_587 = 10'h22f == guard_index ? 64'hf : _GEN_586; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_588 = 10'h230 == guard_index ? 64'h0 : _GEN_587; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_589 = 10'h231 == guard_index ? 64'h1 : _GEN_588; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_590 = 10'h232 == guard_index ? 64'h2 : _GEN_589; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_591 = 10'h233 == guard_index ? 64'h3 : _GEN_590; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_592 = 10'h234 == guard_index ? 64'h4 : _GEN_591; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_593 = 10'h235 == guard_index ? 64'h5 : _GEN_592; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_594 = 10'h236 == guard_index ? 64'h6 : _GEN_593; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_595 = 10'h237 == guard_index ? 64'h7 : _GEN_594; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_596 = 10'h238 == guard_index ? 64'h8 : _GEN_595; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_597 = 10'h239 == guard_index ? 64'h9 : _GEN_596; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_598 = 10'h23a == guard_index ? 64'ha : _GEN_597; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_599 = 10'h23b == guard_index ? 64'hb : _GEN_598; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_600 = 10'h23c == guard_index ? 64'hc : _GEN_599; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_601 = 10'h23d == guard_index ? 64'hd : _GEN_600; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_602 = 10'h23e == guard_index ? 64'he : _GEN_601; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_603 = 10'h23f == guard_index ? 64'hf : _GEN_602; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_604 = 10'h240 == guard_index ? 64'h0 : _GEN_603; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_605 = 10'h241 == guard_index ? 64'h1 : _GEN_604; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_606 = 10'h242 == guard_index ? 64'h2 : _GEN_605; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_607 = 10'h243 == guard_index ? 64'h3 : _GEN_606; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_608 = 10'h244 == guard_index ? 64'h4 : _GEN_607; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_609 = 10'h245 == guard_index ? 64'h5 : _GEN_608; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_610 = 10'h246 == guard_index ? 64'h6 : _GEN_609; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_611 = 10'h247 == guard_index ? 64'h7 : _GEN_610; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_612 = 10'h248 == guard_index ? 64'h8 : _GEN_611; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_613 = 10'h249 == guard_index ? 64'h9 : _GEN_612; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_614 = 10'h24a == guard_index ? 64'ha : _GEN_613; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_615 = 10'h24b == guard_index ? 64'hb : _GEN_614; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_616 = 10'h24c == guard_index ? 64'hc : _GEN_615; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_617 = 10'h24d == guard_index ? 64'hd : _GEN_616; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_618 = 10'h24e == guard_index ? 64'he : _GEN_617; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_619 = 10'h24f == guard_index ? 64'hf : _GEN_618; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_620 = 10'h250 == guard_index ? 64'h0 : _GEN_619; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_621 = 10'h251 == guard_index ? 64'h1 : _GEN_620; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_622 = 10'h252 == guard_index ? 64'h2 : _GEN_621; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_623 = 10'h253 == guard_index ? 64'h3 : _GEN_622; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_624 = 10'h254 == guard_index ? 64'h4 : _GEN_623; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_625 = 10'h255 == guard_index ? 64'h5 : _GEN_624; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_626 = 10'h256 == guard_index ? 64'h6 : _GEN_625; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_627 = 10'h257 == guard_index ? 64'h7 : _GEN_626; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_628 = 10'h258 == guard_index ? 64'h8 : _GEN_627; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_629 = 10'h259 == guard_index ? 64'h9 : _GEN_628; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_630 = 10'h25a == guard_index ? 64'ha : _GEN_629; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_631 = 10'h25b == guard_index ? 64'hb : _GEN_630; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_632 = 10'h25c == guard_index ? 64'hc : _GEN_631; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_633 = 10'h25d == guard_index ? 64'hd : _GEN_632; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_634 = 10'h25e == guard_index ? 64'he : _GEN_633; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_635 = 10'h25f == guard_index ? 64'hf : _GEN_634; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_636 = 10'h260 == guard_index ? 64'h0 : _GEN_635; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_637 = 10'h261 == guard_index ? 64'h1 : _GEN_636; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_638 = 10'h262 == guard_index ? 64'h2 : _GEN_637; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_639 = 10'h263 == guard_index ? 64'h3 : _GEN_638; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_640 = 10'h264 == guard_index ? 64'h4 : _GEN_639; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_641 = 10'h265 == guard_index ? 64'h5 : _GEN_640; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_642 = 10'h266 == guard_index ? 64'h6 : _GEN_641; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_643 = 10'h267 == guard_index ? 64'h7 : _GEN_642; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_644 = 10'h268 == guard_index ? 64'h8 : _GEN_643; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_645 = 10'h269 == guard_index ? 64'h9 : _GEN_644; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_646 = 10'h26a == guard_index ? 64'ha : _GEN_645; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_647 = 10'h26b == guard_index ? 64'hb : _GEN_646; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_648 = 10'h26c == guard_index ? 64'hc : _GEN_647; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_649 = 10'h26d == guard_index ? 64'hd : _GEN_648; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_650 = 10'h26e == guard_index ? 64'he : _GEN_649; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_651 = 10'h26f == guard_index ? 64'hf : _GEN_650; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_652 = 10'h270 == guard_index ? 64'h0 : _GEN_651; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_653 = 10'h271 == guard_index ? 64'h1 : _GEN_652; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_654 = 10'h272 == guard_index ? 64'h2 : _GEN_653; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_655 = 10'h273 == guard_index ? 64'h3 : _GEN_654; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_656 = 10'h274 == guard_index ? 64'h4 : _GEN_655; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_657 = 10'h275 == guard_index ? 64'h5 : _GEN_656; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_658 = 10'h276 == guard_index ? 64'h6 : _GEN_657; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_659 = 10'h277 == guard_index ? 64'h7 : _GEN_658; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_660 = 10'h278 == guard_index ? 64'h8 : _GEN_659; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_661 = 10'h279 == guard_index ? 64'h9 : _GEN_660; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_662 = 10'h27a == guard_index ? 64'ha : _GEN_661; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_663 = 10'h27b == guard_index ? 64'hb : _GEN_662; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_664 = 10'h27c == guard_index ? 64'hc : _GEN_663; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_665 = 10'h27d == guard_index ? 64'hd : _GEN_664; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_666 = 10'h27e == guard_index ? 64'he : _GEN_665; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_667 = 10'h27f == guard_index ? 64'hf : _GEN_666; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_668 = 10'h280 == guard_index ? 64'h0 : _GEN_667; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_669 = 10'h281 == guard_index ? 64'h1 : _GEN_668; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_670 = 10'h282 == guard_index ? 64'h2 : _GEN_669; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_671 = 10'h283 == guard_index ? 64'h3 : _GEN_670; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_672 = 10'h284 == guard_index ? 64'h4 : _GEN_671; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_673 = 10'h285 == guard_index ? 64'h5 : _GEN_672; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_674 = 10'h286 == guard_index ? 64'h6 : _GEN_673; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_675 = 10'h287 == guard_index ? 64'h7 : _GEN_674; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_676 = 10'h288 == guard_index ? 64'h8 : _GEN_675; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_677 = 10'h289 == guard_index ? 64'h9 : _GEN_676; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_678 = 10'h28a == guard_index ? 64'ha : _GEN_677; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_679 = 10'h28b == guard_index ? 64'hb : _GEN_678; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_680 = 10'h28c == guard_index ? 64'hc : _GEN_679; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_681 = 10'h28d == guard_index ? 64'hd : _GEN_680; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_682 = 10'h28e == guard_index ? 64'he : _GEN_681; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_683 = 10'h28f == guard_index ? 64'hf : _GEN_682; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_684 = 10'h290 == guard_index ? 64'h0 : _GEN_683; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_685 = 10'h291 == guard_index ? 64'h1 : _GEN_684; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_686 = 10'h292 == guard_index ? 64'h2 : _GEN_685; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_687 = 10'h293 == guard_index ? 64'h3 : _GEN_686; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_688 = 10'h294 == guard_index ? 64'h4 : _GEN_687; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_689 = 10'h295 == guard_index ? 64'h5 : _GEN_688; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_690 = 10'h296 == guard_index ? 64'h6 : _GEN_689; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_691 = 10'h297 == guard_index ? 64'h7 : _GEN_690; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_692 = 10'h298 == guard_index ? 64'h8 : _GEN_691; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_693 = 10'h299 == guard_index ? 64'h9 : _GEN_692; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_694 = 10'h29a == guard_index ? 64'ha : _GEN_693; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_695 = 10'h29b == guard_index ? 64'hb : _GEN_694; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_696 = 10'h29c == guard_index ? 64'hc : _GEN_695; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_697 = 10'h29d == guard_index ? 64'hd : _GEN_696; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_698 = 10'h29e == guard_index ? 64'he : _GEN_697; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_699 = 10'h29f == guard_index ? 64'hf : _GEN_698; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_700 = 10'h2a0 == guard_index ? 64'h0 : _GEN_699; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_701 = 10'h2a1 == guard_index ? 64'h1 : _GEN_700; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_702 = 10'h2a2 == guard_index ? 64'h2 : _GEN_701; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_703 = 10'h2a3 == guard_index ? 64'h3 : _GEN_702; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_704 = 10'h2a4 == guard_index ? 64'h4 : _GEN_703; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_705 = 10'h2a5 == guard_index ? 64'h5 : _GEN_704; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_706 = 10'h2a6 == guard_index ? 64'h6 : _GEN_705; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_707 = 10'h2a7 == guard_index ? 64'h7 : _GEN_706; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_708 = 10'h2a8 == guard_index ? 64'h8 : _GEN_707; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_709 = 10'h2a9 == guard_index ? 64'h9 : _GEN_708; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_710 = 10'h2aa == guard_index ? 64'ha : _GEN_709; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_711 = 10'h2ab == guard_index ? 64'hb : _GEN_710; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_712 = 10'h2ac == guard_index ? 64'hc : _GEN_711; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_713 = 10'h2ad == guard_index ? 64'hd : _GEN_712; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_714 = 10'h2ae == guard_index ? 64'he : _GEN_713; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_715 = 10'h2af == guard_index ? 64'hf : _GEN_714; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_716 = 10'h2b0 == guard_index ? 64'h0 : _GEN_715; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_717 = 10'h2b1 == guard_index ? 64'h1 : _GEN_716; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_718 = 10'h2b2 == guard_index ? 64'h2 : _GEN_717; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_719 = 10'h2b3 == guard_index ? 64'h3 : _GEN_718; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_720 = 10'h2b4 == guard_index ? 64'h4 : _GEN_719; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_721 = 10'h2b5 == guard_index ? 64'h5 : _GEN_720; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_722 = 10'h2b6 == guard_index ? 64'h6 : _GEN_721; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_723 = 10'h2b7 == guard_index ? 64'h7 : _GEN_722; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_724 = 10'h2b8 == guard_index ? 64'h8 : _GEN_723; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_725 = 10'h2b9 == guard_index ? 64'h9 : _GEN_724; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_726 = 10'h2ba == guard_index ? 64'ha : _GEN_725; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_727 = 10'h2bb == guard_index ? 64'hb : _GEN_726; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_728 = 10'h2bc == guard_index ? 64'hc : _GEN_727; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_729 = 10'h2bd == guard_index ? 64'hd : _GEN_728; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_730 = 10'h2be == guard_index ? 64'he : _GEN_729; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_731 = 10'h2bf == guard_index ? 64'hf : _GEN_730; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_732 = 10'h2c0 == guard_index ? 64'h0 : _GEN_731; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_733 = 10'h2c1 == guard_index ? 64'h1 : _GEN_732; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_734 = 10'h2c2 == guard_index ? 64'h2 : _GEN_733; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_735 = 10'h2c3 == guard_index ? 64'h3 : _GEN_734; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_736 = 10'h2c4 == guard_index ? 64'h4 : _GEN_735; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_737 = 10'h2c5 == guard_index ? 64'h5 : _GEN_736; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_738 = 10'h2c6 == guard_index ? 64'h6 : _GEN_737; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_739 = 10'h2c7 == guard_index ? 64'h7 : _GEN_738; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_740 = 10'h2c8 == guard_index ? 64'h8 : _GEN_739; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_741 = 10'h2c9 == guard_index ? 64'h9 : _GEN_740; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_742 = 10'h2ca == guard_index ? 64'ha : _GEN_741; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_743 = 10'h2cb == guard_index ? 64'hb : _GEN_742; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_744 = 10'h2cc == guard_index ? 64'hc : _GEN_743; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_745 = 10'h2cd == guard_index ? 64'hd : _GEN_744; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_746 = 10'h2ce == guard_index ? 64'he : _GEN_745; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_747 = 10'h2cf == guard_index ? 64'hf : _GEN_746; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_748 = 10'h2d0 == guard_index ? 64'h0 : _GEN_747; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_749 = 10'h2d1 == guard_index ? 64'h1 : _GEN_748; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_750 = 10'h2d2 == guard_index ? 64'h2 : _GEN_749; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_751 = 10'h2d3 == guard_index ? 64'h3 : _GEN_750; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_752 = 10'h2d4 == guard_index ? 64'h4 : _GEN_751; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_753 = 10'h2d5 == guard_index ? 64'h5 : _GEN_752; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_754 = 10'h2d6 == guard_index ? 64'h6 : _GEN_753; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_755 = 10'h2d7 == guard_index ? 64'h7 : _GEN_754; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_756 = 10'h2d8 == guard_index ? 64'h8 : _GEN_755; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_757 = 10'h2d9 == guard_index ? 64'h9 : _GEN_756; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_758 = 10'h2da == guard_index ? 64'ha : _GEN_757; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_759 = 10'h2db == guard_index ? 64'hb : _GEN_758; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_760 = 10'h2dc == guard_index ? 64'hc : _GEN_759; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_761 = 10'h2dd == guard_index ? 64'hd : _GEN_760; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_762 = 10'h2de == guard_index ? 64'he : _GEN_761; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_763 = 10'h2df == guard_index ? 64'hf : _GEN_762; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_764 = 10'h2e0 == guard_index ? 64'h0 : _GEN_763; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_765 = 10'h2e1 == guard_index ? 64'h1 : _GEN_764; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_766 = 10'h2e2 == guard_index ? 64'h2 : _GEN_765; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_767 = 10'h2e3 == guard_index ? 64'h3 : _GEN_766; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_768 = 10'h2e4 == guard_index ? 64'h4 : _GEN_767; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_769 = 10'h2e5 == guard_index ? 64'h5 : _GEN_768; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_770 = 10'h2e6 == guard_index ? 64'h6 : _GEN_769; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_771 = 10'h2e7 == guard_index ? 64'h7 : _GEN_770; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_772 = 10'h2e8 == guard_index ? 64'h8 : _GEN_771; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_773 = 10'h2e9 == guard_index ? 64'h9 : _GEN_772; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_774 = 10'h2ea == guard_index ? 64'ha : _GEN_773; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_775 = 10'h2eb == guard_index ? 64'hb : _GEN_774; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_776 = 10'h2ec == guard_index ? 64'hc : _GEN_775; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_777 = 10'h2ed == guard_index ? 64'hd : _GEN_776; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_778 = 10'h2ee == guard_index ? 64'he : _GEN_777; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_779 = 10'h2ef == guard_index ? 64'hf : _GEN_778; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_780 = 10'h2f0 == guard_index ? 64'h0 : _GEN_779; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_781 = 10'h2f1 == guard_index ? 64'h1 : _GEN_780; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_782 = 10'h2f2 == guard_index ? 64'h2 : _GEN_781; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_783 = 10'h2f3 == guard_index ? 64'h3 : _GEN_782; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_784 = 10'h2f4 == guard_index ? 64'h4 : _GEN_783; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_785 = 10'h2f5 == guard_index ? 64'h5 : _GEN_784; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_786 = 10'h2f6 == guard_index ? 64'h6 : _GEN_785; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_787 = 10'h2f7 == guard_index ? 64'h7 : _GEN_786; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_788 = 10'h2f8 == guard_index ? 64'h8 : _GEN_787; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_789 = 10'h2f9 == guard_index ? 64'h9 : _GEN_788; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_790 = 10'h2fa == guard_index ? 64'ha : _GEN_789; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_791 = 10'h2fb == guard_index ? 64'hb : _GEN_790; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_792 = 10'h2fc == guard_index ? 64'hc : _GEN_791; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_793 = 10'h2fd == guard_index ? 64'hd : _GEN_792; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_794 = 10'h2fe == guard_index ? 64'he : _GEN_793; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_795 = 10'h2ff == guard_index ? 64'hf : _GEN_794; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_796 = 10'h300 == guard_index ? 64'h0 : _GEN_795; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_797 = 10'h301 == guard_index ? 64'h1 : _GEN_796; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_798 = 10'h302 == guard_index ? 64'h2 : _GEN_797; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_799 = 10'h303 == guard_index ? 64'h3 : _GEN_798; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_800 = 10'h304 == guard_index ? 64'h4 : _GEN_799; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_801 = 10'h305 == guard_index ? 64'h5 : _GEN_800; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_802 = 10'h306 == guard_index ? 64'h6 : _GEN_801; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_803 = 10'h307 == guard_index ? 64'h7 : _GEN_802; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_804 = 10'h308 == guard_index ? 64'h8 : _GEN_803; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_805 = 10'h309 == guard_index ? 64'h9 : _GEN_804; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_806 = 10'h30a == guard_index ? 64'ha : _GEN_805; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_807 = 10'h30b == guard_index ? 64'hb : _GEN_806; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_808 = 10'h30c == guard_index ? 64'hc : _GEN_807; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_809 = 10'h30d == guard_index ? 64'hd : _GEN_808; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_810 = 10'h30e == guard_index ? 64'he : _GEN_809; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_811 = 10'h30f == guard_index ? 64'hf : _GEN_810; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_812 = 10'h310 == guard_index ? 64'h0 : _GEN_811; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_813 = 10'h311 == guard_index ? 64'h1 : _GEN_812; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_814 = 10'h312 == guard_index ? 64'h2 : _GEN_813; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_815 = 10'h313 == guard_index ? 64'h3 : _GEN_814; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_816 = 10'h314 == guard_index ? 64'h4 : _GEN_815; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_817 = 10'h315 == guard_index ? 64'h5 : _GEN_816; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_818 = 10'h316 == guard_index ? 64'h6 : _GEN_817; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_819 = 10'h317 == guard_index ? 64'h7 : _GEN_818; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_820 = 10'h318 == guard_index ? 64'h8 : _GEN_819; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_821 = 10'h319 == guard_index ? 64'h9 : _GEN_820; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_822 = 10'h31a == guard_index ? 64'ha : _GEN_821; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_823 = 10'h31b == guard_index ? 64'hb : _GEN_822; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_824 = 10'h31c == guard_index ? 64'hc : _GEN_823; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_825 = 10'h31d == guard_index ? 64'hd : _GEN_824; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_826 = 10'h31e == guard_index ? 64'he : _GEN_825; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_827 = 10'h31f == guard_index ? 64'hf : _GEN_826; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_828 = 10'h320 == guard_index ? 64'h0 : _GEN_827; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_829 = 10'h321 == guard_index ? 64'h1 : _GEN_828; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_830 = 10'h322 == guard_index ? 64'h2 : _GEN_829; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_831 = 10'h323 == guard_index ? 64'h3 : _GEN_830; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_832 = 10'h324 == guard_index ? 64'h4 : _GEN_831; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_833 = 10'h325 == guard_index ? 64'h5 : _GEN_832; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_834 = 10'h326 == guard_index ? 64'h6 : _GEN_833; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_835 = 10'h327 == guard_index ? 64'h7 : _GEN_834; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_836 = 10'h328 == guard_index ? 64'h8 : _GEN_835; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_837 = 10'h329 == guard_index ? 64'h9 : _GEN_836; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_838 = 10'h32a == guard_index ? 64'ha : _GEN_837; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_839 = 10'h32b == guard_index ? 64'hb : _GEN_838; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_840 = 10'h32c == guard_index ? 64'hc : _GEN_839; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_841 = 10'h32d == guard_index ? 64'hd : _GEN_840; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_842 = 10'h32e == guard_index ? 64'he : _GEN_841; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_843 = 10'h32f == guard_index ? 64'hf : _GEN_842; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_844 = 10'h330 == guard_index ? 64'h0 : _GEN_843; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_845 = 10'h331 == guard_index ? 64'h1 : _GEN_844; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_846 = 10'h332 == guard_index ? 64'h2 : _GEN_845; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_847 = 10'h333 == guard_index ? 64'h3 : _GEN_846; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_848 = 10'h334 == guard_index ? 64'h4 : _GEN_847; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_849 = 10'h335 == guard_index ? 64'h5 : _GEN_848; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_850 = 10'h336 == guard_index ? 64'h6 : _GEN_849; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_851 = 10'h337 == guard_index ? 64'h7 : _GEN_850; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_852 = 10'h338 == guard_index ? 64'h8 : _GEN_851; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_853 = 10'h339 == guard_index ? 64'h9 : _GEN_852; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_854 = 10'h33a == guard_index ? 64'ha : _GEN_853; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_855 = 10'h33b == guard_index ? 64'hb : _GEN_854; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_856 = 10'h33c == guard_index ? 64'hc : _GEN_855; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_857 = 10'h33d == guard_index ? 64'hd : _GEN_856; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_858 = 10'h33e == guard_index ? 64'he : _GEN_857; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_859 = 10'h33f == guard_index ? 64'hf : _GEN_858; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_860 = 10'h340 == guard_index ? 64'h0 : _GEN_859; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_861 = 10'h341 == guard_index ? 64'h1 : _GEN_860; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_862 = 10'h342 == guard_index ? 64'h2 : _GEN_861; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_863 = 10'h343 == guard_index ? 64'h3 : _GEN_862; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_864 = 10'h344 == guard_index ? 64'h4 : _GEN_863; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_865 = 10'h345 == guard_index ? 64'h5 : _GEN_864; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_866 = 10'h346 == guard_index ? 64'h6 : _GEN_865; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_867 = 10'h347 == guard_index ? 64'h7 : _GEN_866; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_868 = 10'h348 == guard_index ? 64'h8 : _GEN_867; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_869 = 10'h349 == guard_index ? 64'h9 : _GEN_868; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_870 = 10'h34a == guard_index ? 64'ha : _GEN_869; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_871 = 10'h34b == guard_index ? 64'hb : _GEN_870; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_872 = 10'h34c == guard_index ? 64'hc : _GEN_871; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_873 = 10'h34d == guard_index ? 64'hd : _GEN_872; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_874 = 10'h34e == guard_index ? 64'he : _GEN_873; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_875 = 10'h34f == guard_index ? 64'hf : _GEN_874; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_876 = 10'h350 == guard_index ? 64'h0 : _GEN_875; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_877 = 10'h351 == guard_index ? 64'h1 : _GEN_876; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_878 = 10'h352 == guard_index ? 64'h2 : _GEN_877; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_879 = 10'h353 == guard_index ? 64'h3 : _GEN_878; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_880 = 10'h354 == guard_index ? 64'h4 : _GEN_879; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_881 = 10'h355 == guard_index ? 64'h5 : _GEN_880; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_882 = 10'h356 == guard_index ? 64'h6 : _GEN_881; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_883 = 10'h357 == guard_index ? 64'h7 : _GEN_882; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_884 = 10'h358 == guard_index ? 64'h8 : _GEN_883; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_885 = 10'h359 == guard_index ? 64'h9 : _GEN_884; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_886 = 10'h35a == guard_index ? 64'ha : _GEN_885; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_887 = 10'h35b == guard_index ? 64'hb : _GEN_886; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_888 = 10'h35c == guard_index ? 64'hc : _GEN_887; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_889 = 10'h35d == guard_index ? 64'hd : _GEN_888; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_890 = 10'h35e == guard_index ? 64'he : _GEN_889; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_891 = 10'h35f == guard_index ? 64'hf : _GEN_890; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_892 = 10'h360 == guard_index ? 64'h0 : _GEN_891; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_893 = 10'h361 == guard_index ? 64'h1 : _GEN_892; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_894 = 10'h362 == guard_index ? 64'h2 : _GEN_893; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_895 = 10'h363 == guard_index ? 64'h3 : _GEN_894; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_896 = 10'h364 == guard_index ? 64'h4 : _GEN_895; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_897 = 10'h365 == guard_index ? 64'h5 : _GEN_896; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_898 = 10'h366 == guard_index ? 64'h6 : _GEN_897; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_899 = 10'h367 == guard_index ? 64'h7 : _GEN_898; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_900 = 10'h368 == guard_index ? 64'h8 : _GEN_899; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_901 = 10'h369 == guard_index ? 64'h9 : _GEN_900; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_902 = 10'h36a == guard_index ? 64'ha : _GEN_901; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_903 = 10'h36b == guard_index ? 64'hb : _GEN_902; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_904 = 10'h36c == guard_index ? 64'hc : _GEN_903; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_905 = 10'h36d == guard_index ? 64'hd : _GEN_904; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_906 = 10'h36e == guard_index ? 64'he : _GEN_905; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_907 = 10'h36f == guard_index ? 64'hf : _GEN_906; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_908 = 10'h370 == guard_index ? 64'h0 : _GEN_907; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_909 = 10'h371 == guard_index ? 64'h1 : _GEN_908; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_910 = 10'h372 == guard_index ? 64'h2 : _GEN_909; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_911 = 10'h373 == guard_index ? 64'h3 : _GEN_910; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_912 = 10'h374 == guard_index ? 64'h4 : _GEN_911; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_913 = 10'h375 == guard_index ? 64'h5 : _GEN_912; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_914 = 10'h376 == guard_index ? 64'h6 : _GEN_913; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_915 = 10'h377 == guard_index ? 64'h7 : _GEN_914; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_916 = 10'h378 == guard_index ? 64'h8 : _GEN_915; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_917 = 10'h379 == guard_index ? 64'h9 : _GEN_916; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_918 = 10'h37a == guard_index ? 64'ha : _GEN_917; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_919 = 10'h37b == guard_index ? 64'hb : _GEN_918; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_920 = 10'h37c == guard_index ? 64'hc : _GEN_919; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_921 = 10'h37d == guard_index ? 64'hd : _GEN_920; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_922 = 10'h37e == guard_index ? 64'he : _GEN_921; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_923 = 10'h37f == guard_index ? 64'hf : _GEN_922; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_924 = 10'h380 == guard_index ? 64'h0 : _GEN_923; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_925 = 10'h381 == guard_index ? 64'h1 : _GEN_924; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_926 = 10'h382 == guard_index ? 64'h2 : _GEN_925; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_927 = 10'h383 == guard_index ? 64'h3 : _GEN_926; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_928 = 10'h384 == guard_index ? 64'h4 : _GEN_927; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_929 = 10'h385 == guard_index ? 64'h5 : _GEN_928; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_930 = 10'h386 == guard_index ? 64'h6 : _GEN_929; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_931 = 10'h387 == guard_index ? 64'h7 : _GEN_930; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_932 = 10'h388 == guard_index ? 64'h8 : _GEN_931; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_933 = 10'h389 == guard_index ? 64'h9 : _GEN_932; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_934 = 10'h38a == guard_index ? 64'ha : _GEN_933; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_935 = 10'h38b == guard_index ? 64'hb : _GEN_934; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_936 = 10'h38c == guard_index ? 64'hc : _GEN_935; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_937 = 10'h38d == guard_index ? 64'hd : _GEN_936; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_938 = 10'h38e == guard_index ? 64'he : _GEN_937; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_939 = 10'h38f == guard_index ? 64'hf : _GEN_938; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_940 = 10'h390 == guard_index ? 64'h0 : _GEN_939; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_941 = 10'h391 == guard_index ? 64'h1 : _GEN_940; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_942 = 10'h392 == guard_index ? 64'h2 : _GEN_941; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_943 = 10'h393 == guard_index ? 64'h3 : _GEN_942; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_944 = 10'h394 == guard_index ? 64'h4 : _GEN_943; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_945 = 10'h395 == guard_index ? 64'h5 : _GEN_944; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_946 = 10'h396 == guard_index ? 64'h6 : _GEN_945; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_947 = 10'h397 == guard_index ? 64'h7 : _GEN_946; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_948 = 10'h398 == guard_index ? 64'h8 : _GEN_947; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_949 = 10'h399 == guard_index ? 64'h9 : _GEN_948; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_950 = 10'h39a == guard_index ? 64'ha : _GEN_949; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_951 = 10'h39b == guard_index ? 64'hb : _GEN_950; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_952 = 10'h39c == guard_index ? 64'hc : _GEN_951; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_953 = 10'h39d == guard_index ? 64'hd : _GEN_952; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_954 = 10'h39e == guard_index ? 64'he : _GEN_953; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_955 = 10'h39f == guard_index ? 64'hf : _GEN_954; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_956 = 10'h3a0 == guard_index ? 64'h0 : _GEN_955; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_957 = 10'h3a1 == guard_index ? 64'h1 : _GEN_956; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_958 = 10'h3a2 == guard_index ? 64'h2 : _GEN_957; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_959 = 10'h3a3 == guard_index ? 64'h3 : _GEN_958; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_960 = 10'h3a4 == guard_index ? 64'h4 : _GEN_959; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_961 = 10'h3a5 == guard_index ? 64'h5 : _GEN_960; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_962 = 10'h3a6 == guard_index ? 64'h6 : _GEN_961; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_963 = 10'h3a7 == guard_index ? 64'h7 : _GEN_962; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_964 = 10'h3a8 == guard_index ? 64'h8 : _GEN_963; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_965 = 10'h3a9 == guard_index ? 64'h9 : _GEN_964; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_966 = 10'h3aa == guard_index ? 64'ha : _GEN_965; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_967 = 10'h3ab == guard_index ? 64'hb : _GEN_966; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_968 = 10'h3ac == guard_index ? 64'hc : _GEN_967; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_969 = 10'h3ad == guard_index ? 64'hd : _GEN_968; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_970 = 10'h3ae == guard_index ? 64'he : _GEN_969; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_971 = 10'h3af == guard_index ? 64'hf : _GEN_970; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_972 = 10'h3b0 == guard_index ? 64'h0 : _GEN_971; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_973 = 10'h3b1 == guard_index ? 64'h1 : _GEN_972; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_974 = 10'h3b2 == guard_index ? 64'h2 : _GEN_973; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_975 = 10'h3b3 == guard_index ? 64'h3 : _GEN_974; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_976 = 10'h3b4 == guard_index ? 64'h4 : _GEN_975; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_977 = 10'h3b5 == guard_index ? 64'h5 : _GEN_976; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_978 = 10'h3b6 == guard_index ? 64'h6 : _GEN_977; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_979 = 10'h3b7 == guard_index ? 64'h7 : _GEN_978; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_980 = 10'h3b8 == guard_index ? 64'h8 : _GEN_979; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_981 = 10'h3b9 == guard_index ? 64'h9 : _GEN_980; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_982 = 10'h3ba == guard_index ? 64'ha : _GEN_981; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_983 = 10'h3bb == guard_index ? 64'hb : _GEN_982; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_984 = 10'h3bc == guard_index ? 64'hc : _GEN_983; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_985 = 10'h3bd == guard_index ? 64'hd : _GEN_984; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_986 = 10'h3be == guard_index ? 64'he : _GEN_985; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_987 = 10'h3bf == guard_index ? 64'hf : _GEN_986; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_988 = 10'h3c0 == guard_index ? 64'h0 : _GEN_987; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_989 = 10'h3c1 == guard_index ? 64'h1 : _GEN_988; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_990 = 10'h3c2 == guard_index ? 64'h2 : _GEN_989; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_991 = 10'h3c3 == guard_index ? 64'h3 : _GEN_990; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_992 = 10'h3c4 == guard_index ? 64'h4 : _GEN_991; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_993 = 10'h3c5 == guard_index ? 64'h5 : _GEN_992; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_994 = 10'h3c6 == guard_index ? 64'h6 : _GEN_993; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_995 = 10'h3c7 == guard_index ? 64'h7 : _GEN_994; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_996 = 10'h3c8 == guard_index ? 64'h8 : _GEN_995; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_997 = 10'h3c9 == guard_index ? 64'h9 : _GEN_996; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_998 = 10'h3ca == guard_index ? 64'ha : _GEN_997; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_999 = 10'h3cb == guard_index ? 64'hb : _GEN_998; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1000 = 10'h3cc == guard_index ? 64'hc : _GEN_999; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1001 = 10'h3cd == guard_index ? 64'hd : _GEN_1000; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1002 = 10'h3ce == guard_index ? 64'he : _GEN_1001; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1003 = 10'h3cf == guard_index ? 64'hf : _GEN_1002; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1004 = 10'h3d0 == guard_index ? 64'h0 : _GEN_1003; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1005 = 10'h3d1 == guard_index ? 64'h1 : _GEN_1004; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1006 = 10'h3d2 == guard_index ? 64'h2 : _GEN_1005; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1007 = 10'h3d3 == guard_index ? 64'h3 : _GEN_1006; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1008 = 10'h3d4 == guard_index ? 64'h4 : _GEN_1007; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1009 = 10'h3d5 == guard_index ? 64'h5 : _GEN_1008; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1010 = 10'h3d6 == guard_index ? 64'h6 : _GEN_1009; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1011 = 10'h3d7 == guard_index ? 64'h7 : _GEN_1010; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1012 = 10'h3d8 == guard_index ? 64'h8 : _GEN_1011; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1013 = 10'h3d9 == guard_index ? 64'h9 : _GEN_1012; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1014 = 10'h3da == guard_index ? 64'ha : _GEN_1013; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1015 = 10'h3db == guard_index ? 64'hb : _GEN_1014; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1016 = 10'h3dc == guard_index ? 64'hc : _GEN_1015; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1017 = 10'h3dd == guard_index ? 64'hd : _GEN_1016; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1018 = 10'h3de == guard_index ? 64'he : _GEN_1017; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1019 = 10'h3df == guard_index ? 64'hf : _GEN_1018; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1020 = 10'h3e0 == guard_index ? 64'h0 : _GEN_1019; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1021 = 10'h3e1 == guard_index ? 64'h1 : _GEN_1020; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1022 = 10'h3e2 == guard_index ? 64'h2 : _GEN_1021; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1023 = 10'h3e3 == guard_index ? 64'h3 : _GEN_1022; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1024 = 10'h3e4 == guard_index ? 64'h4 : _GEN_1023; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1025 = 10'h3e5 == guard_index ? 64'h5 : _GEN_1024; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1026 = 10'h3e6 == guard_index ? 64'h6 : _GEN_1025; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1027 = 10'h3e7 == guard_index ? 64'h7 : _GEN_1026; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1028 = 10'h3e8 == guard_index ? 64'h8 : _GEN_1027; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1029 = 10'h3e9 == guard_index ? 64'h9 : _GEN_1028; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1030 = 10'h3ea == guard_index ? 64'ha : _GEN_1029; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1031 = 10'h3eb == guard_index ? 64'hb : _GEN_1030; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1032 = 10'h3ec == guard_index ? 64'hc : _GEN_1031; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1033 = 10'h3ed == guard_index ? 64'hd : _GEN_1032; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1034 = 10'h3ee == guard_index ? 64'he : _GEN_1033; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1035 = 10'h3ef == guard_index ? 64'hf : _GEN_1034; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1036 = 10'h3f0 == guard_index ? 64'h0 : _GEN_1035; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1037 = 10'h3f1 == guard_index ? 64'h1 : _GEN_1036; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1038 = 10'h3f2 == guard_index ? 64'h2 : _GEN_1037; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1039 = 10'h3f3 == guard_index ? 64'h3 : _GEN_1038; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1040 = 10'h3f4 == guard_index ? 64'h4 : _GEN_1039; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1041 = 10'h3f5 == guard_index ? 64'h5 : _GEN_1040; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1042 = 10'h3f6 == guard_index ? 64'h6 : _GEN_1041; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1043 = 10'h3f7 == guard_index ? 64'h7 : _GEN_1042; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1044 = 10'h3f8 == guard_index ? 64'h8 : _GEN_1043; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1045 = 10'h3f9 == guard_index ? 64'h9 : _GEN_1044; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1046 = 10'h3fa == guard_index ? 64'ha : _GEN_1045; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1047 = 10'h3fb == guard_index ? 64'hb : _GEN_1046; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1048 = 10'h3fc == guard_index ? 64'hc : _GEN_1047; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1049 = 10'h3fd == guard_index ? 64'hd : _GEN_1048; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1050 = 10'h3fe == guard_index ? 64'he : _GEN_1049; // @[PhiNode.scala 336:38]
  wire [63:0] _GEN_1051 = 10'h3ff == guard_index ? 64'hf : _GEN_1050; // @[PhiNode.scala 336:38]
  wire  _T_45 = _GEN_27 != _GEN_1051; // @[PhiNode.scala 336:38]
  wire  _T_34 = _T_43 & enable_R_control; // @[PhiNode.scala 290:38]
  wire  _T_35 = state == 2'h0; // @[PhiNode.scala 290:67]
  wire  _T_36 = _T_34 & _T_35; // @[PhiNode.scala 290:58]
  wire [9:0] _T_40 = guard_index + 10'h1; // @[Counter.scala 39:22]
  wire [4:0] _GEN_26 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 312:12]
  wire  _T_47 = ~reset; // @[PhiNode.scala 341:23]
  wire [4:0] _GEN_1062 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 350:19]
  wire  _GEN_1067 = _T_43 | _GEN_17; // @[PhiNode.scala 327:66]
  wire  _GEN_1068 = _T_43 | _GEN_19; // @[PhiNode.scala 327:66]
  wire  _T_52 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 364:31]
  wire  _T_57 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_1107 = _T_57 ? 64'h0 : _GEN_27; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_1148 = _T_52 ? _GEN_27 : _GEN_1107; // @[Conditional.scala 39:67]
  wire  _GEN_1181 = _T_41 & _T_43; // @[PhiNode.scala 341:23]
  wire  _GEN_1182 = _GEN_1181 & enable_R_control; // @[PhiNode.scala 341:23]
  wire  _GEN_1183 = _GEN_1182 & _T_45; // @[PhiNode.scala 341:23]
  wire  _GEN_1187 = ~enable_R_control; // @[PhiNode.scala 357:19]
  wire  _GEN_1188 = _GEN_1181 & _GEN_1187; // @[PhiNode.scala 357:19]
  assign io_enable_ready = ~enable_valid_R; // @[PhiNode.scala 245:19]
  assign io_InData_0_ready = ~in_data_valid_R_0; // @[PhiNode.scala 253:24]
  assign io_InData_1_ready = ~in_data_valid_R_1; // @[PhiNode.scala 253:24]
  assign io_Mask_ready = ~mask_valid_R; // @[PhiNode.scala 238:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 322:21]
  assign io_Out_0_bits_data = _T_41 ? _GEN_27 : _GEN_1148; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 322:21]
  assign io_Out_1_bits_data = _T_41 ? _GEN_27 : _GEN_1148; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[4:0];
  _RAND_3 = {2{`RANDOM}};
  in_data_R_1_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_R_control = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  enable_valid_R = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mask_R = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  mask_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fire_R_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  guard_index = _RAND_15[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else if (_T_41) begin
      if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        in_data_R_0_taskID <= 5'h0;
      end else if (_T_14) begin
        in_data_R_0_taskID <= io_InData_0_bits_taskID;
      end
    end else if (_T_14) begin
      in_data_R_0_taskID <= io_InData_0_bits_taskID;
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else if (_T_41) begin
      if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        in_data_R_1_taskID <= 5'h0;
      end else if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        in_data_R_1_taskID <= 5'h0;
      end else if (_T_16) begin
        in_data_R_1_taskID <= io_InData_1_bits_taskID;
      end
    end else if (_T_16) begin
      in_data_R_1_taskID <= io_InData_1_bits_taskID;
    end
    if (reset) begin
      in_data_R_1_data <= 64'h0;
    end else if (_T_41) begin
      if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_16) begin
      in_data_R_1_data <= io_InData_1_bits_data;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_41) begin
      in_data_valid_R_0 <= _GEN_11;
    end else if (_T_52) begin
      if (_T_53) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_11;
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else if (_T_41) begin
      in_data_valid_R_1 <= _GEN_15;
    end else if (_T_52) begin
      if (_T_53) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else begin
      in_data_valid_R_1 <= _GEN_15;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_41) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_41) begin
      enable_valid_R <= _GEN_7;
    end else if (_T_52) begin
      if (_T_53) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else begin
      enable_valid_R <= _GEN_7;
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else if (_T_41) begin
      if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_10) begin
      mask_R <= io_Mask_bits;
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else if (_T_41) begin
      mask_valid_R <= _GEN_3;
    end else if (_T_52) begin
      if (_T_53) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else begin
      mask_valid_R <= _GEN_3;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_41) begin
      if (_T_43) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_52) begin
      if (_T_53) begin
        state <= 2'h0;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_41) begin
      out_valid_R_0 <= _GEN_1067;
    end else if (_T_20) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_41) begin
      out_valid_R_1 <= _GEN_1068;
    end else if (_T_21) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else if (_T_41) begin
      fire_R_0 <= _GEN_16;
    end else if (_T_52) begin
      if (_T_53) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else begin
      fire_R_0 <= _GEN_16;
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else if (_T_41) begin
      fire_R_1 <= _GEN_18;
    end else if (_T_52) begin
      if (_T_53) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else if (_T_57) begin
      if (_T_53) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else begin
      fire_R_1 <= _GEN_18;
    end
    if (reset) begin
      guard_index <= 10'h0;
    end else if (_T_36) begin
      guard_index <= _T_40;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1183 & _T_47) begin
          $fwrite(32'h80000002,"[DEBUG] [Bbgemm] [TID->%d] [PHI] phiindvars_iv785 Produced value: %d, correct value: %d\n",_GEN_26,_GEN_27,_GEN_1051); // @[PhiNode.scala 341:23]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1182 & _T_47) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv785] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_1062,enable_R_control,_GEN_27,cycleCount); // @[PhiNode.scala 350:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1188 & _T_47) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv785] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_1062,enable_R_control,_GEN_27,cycleCount); // @[PhiNode.scala 357:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU(
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out
);
  wire [524350:0] _GEN_0 = {{524287'd0}, io_in1}; // @[Alu.scala 183:38]
  wire [524350:0] _T_10 = _GEN_0 << io_in2[18:0]; // @[Alu.scala 183:38]
  assign io_out = _T_10[63:0]; // @[Alu.scala 235:10]
endmodule
module ComputeNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h4;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_6] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: shl] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_3(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  state; // @[BranchNode.scala 588:22]
  wire  _T_11 = ~state; // @[Conditional.scala 37:30]
  wire  _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_16 = ~reset; // @[BranchNode.scala 616:17]
  wire  _GEN_8 = enable_valid_R | state; // @[BranchNode.scala 611:46]
  wire  _GEN_10 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 611:46]
  wire  _T_18 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_19 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_20 = _T_18 | _T_19; // @[HandShaking.scala 725:29]
  wire  _GEN_31 = _T_11 & enable_valid_R; // @[BranchNode.scala 616:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = _T_11 ? _GEN_10 : out_valid_R_0; // @[HandShaking.scala 630:21 BranchNode.scala 614:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 607:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 607:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_control <= 1'h0;
      end else if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_20) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (enable_valid_R) begin
        out_valid_R_0 <= _T_14;
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_11) begin
      state <= _GEN_8;
    end else if (state) begin
      if (_T_20) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [UBR] [br_7] [Out: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,cycleCount); // @[BranchNode.scala 616:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [63:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [63:0] io_Out_2_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] in_data_R_1_data; // @[PhiNode.scala 203:26]
  reg  in_data_valid_R_0; // @[PhiNode.scala 204:32]
  reg  in_data_valid_R_1; // @[PhiNode.scala 204:32]
  reg  enable_R_control; // @[PhiNode.scala 207:25]
  reg  enable_valid_R; // @[PhiNode.scala 208:31]
  reg [1:0] mask_R; // @[PhiNode.scala 211:23]
  reg  mask_valid_R; // @[PhiNode.scala 212:29]
  reg [1:0] state; // @[PhiNode.scala 216:22]
  reg  out_valid_R_0; // @[PhiNode.scala 219:49]
  reg  out_valid_R_1; // @[PhiNode.scala 219:49]
  reg  out_valid_R_2; // @[PhiNode.scala 219:49]
  reg  fire_R_0; // @[PhiNode.scala 221:44]
  reg  fire_R_1; // @[PhiNode.scala 221:44]
  reg  fire_R_2; // @[PhiNode.scala 221:44]
  wire  _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_10 | mask_valid_R; // @[PhiNode.scala 239:24]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_12 | enable_valid_R; // @[PhiNode.scala 246:26]
  wire  _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 254:29]
  wire  _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 254:29]
  wire [1:0] _T_19 = {mask_R[0],mask_R[1]}; // @[Cat.scala 29:58]
  wire  sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  wire  _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_16 = _T_20 | fire_R_0; // @[PhiNode.scala 276:26]
  wire  _GEN_17 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 276:26]
  wire  _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = _T_21 | fire_R_1; // @[PhiNode.scala 276:26]
  wire  _GEN_19 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 276:26]
  wire  _T_22 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_20 = _T_22 | fire_R_2; // @[PhiNode.scala 276:26]
  wire  _GEN_21 = _T_22 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 276:26]
  wire  fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 283:74]
  wire  fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 283:74]
  wire  fire_mask_2 = fire_R_2 | _T_22; // @[PhiNode.scala 283:74]
  wire [63:0] _GEN_28 = sel ? in_data_R_1_data : 64'h0; // @[PhiNode.scala 312:12]
  wire  _T_31 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 286:30]
  wire  _T_32 = enable_valid_R & _T_31; // @[PhiNode.scala 290:20]
  wire  _T_37 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_42 = ~reset; // @[PhiNode.scala 350:19]
  wire [4:0] _GEN_37 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 350:19]
  wire  _GEN_40 = _T_32 | _GEN_17; // @[PhiNode.scala 327:66]
  wire  _GEN_41 = _T_32 | _GEN_19; // @[PhiNode.scala 327:66]
  wire  _GEN_42 = _T_32 | _GEN_21; // @[PhiNode.scala 327:66]
  wire  _T_45 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_46 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 364:31]
  wire  _T_47 = _T_46 & fire_mask_2; // @[PhiNode.scala 364:31]
  wire  _T_51 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_81 = _T_51 ? 64'h0 : _GEN_28; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_127 = _T_45 ? _GEN_28 : _GEN_81; // @[Conditional.scala 39:67]
  wire  _GEN_167 = _T_37 & _T_32; // @[PhiNode.scala 350:19]
  wire  _GEN_168 = _GEN_167 & enable_R_control; // @[PhiNode.scala 350:19]
  wire  _GEN_170 = ~enable_R_control; // @[PhiNode.scala 357:19]
  wire  _GEN_171 = _GEN_167 & _GEN_170; // @[PhiNode.scala 357:19]
  assign io_enable_ready = ~enable_valid_R; // @[PhiNode.scala 245:19]
  assign io_InData_0_ready = ~in_data_valid_R_0; // @[PhiNode.scala 253:24]
  assign io_InData_1_ready = ~in_data_valid_R_1; // @[PhiNode.scala 253:24]
  assign io_Mask_ready = ~mask_valid_R; // @[PhiNode.scala 238:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 322:21]
  assign io_Out_0_bits_data = _T_37 ? _GEN_28 : _GEN_127; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 322:21]
  assign io_Out_1_bits_data = _T_37 ? _GEN_28 : _GEN_127; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 322:21]
  assign io_Out_2_bits_data = _T_37 ? _GEN_28 : _GEN_127; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {2{`RANDOM}};
  in_data_R_1_data = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_R_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fire_R_2 = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_1_data <= 64'h0;
    end else if (_T_37) begin
      if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_45) begin
      if (_T_47) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_16) begin
      in_data_R_1_data <= io_InData_1_bits_data;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      in_data_valid_R_0 <= _GEN_11;
    end else if (_T_45) begin
      if (_T_47) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_11;
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else if (_T_37) begin
      in_data_valid_R_1 <= _GEN_15;
    end else if (_T_45) begin
      if (_T_47) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else begin
      in_data_valid_R_1 <= _GEN_15;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_37) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_45) begin
      if (_T_47) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_37) begin
      enable_valid_R <= _GEN_7;
    end else if (_T_45) begin
      if (_T_47) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else begin
      enable_valid_R <= _GEN_7;
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else if (_T_37) begin
      if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_45) begin
      if (_T_47) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_10) begin
      mask_R <= io_Mask_bits;
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else if (_T_37) begin
      mask_valid_R <= _GEN_3;
    end else if (_T_45) begin
      if (_T_47) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else begin
      mask_valid_R <= _GEN_3;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_37) begin
      if (_T_32) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_45) begin
      if (_T_47) begin
        state <= 2'h0;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_0 <= _GEN_40;
    end else if (_T_20) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_1 <= _GEN_41;
    end else if (_T_21) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_2 <= _GEN_42;
    end else if (_T_22) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else if (_T_37) begin
      fire_R_0 <= _GEN_16;
    end else if (_T_45) begin
      if (_T_47) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else begin
      fire_R_0 <= _GEN_16;
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else if (_T_37) begin
      fire_R_1 <= _GEN_18;
    end else if (_T_45) begin
      if (_T_47) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else begin
      fire_R_1 <= _GEN_18;
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else if (_T_37) begin
      fire_R_2 <= _GEN_20;
    end else if (_T_45) begin
      if (_T_47) begin
        fire_R_2 <= 1'h0;
      end else begin
        fire_R_2 <= _GEN_20;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        fire_R_2 <= 1'h0;
      end else begin
        fire_R_2 <= _GEN_20;
      end
    end else begin
      fire_R_2 <= _GEN_20;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_168 & _T_42) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv718] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_37,enable_R_control,_GEN_28,cycleCount); // @[PhiNode.scala 350:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_42) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv718] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_37,enable_R_control,_GEN_28,cycleCount); // @[PhiNode.scala 357:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_1(
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out
);
  assign io_out = io_in1 + io_in2; // @[Alu.scala 235:10]
endmodule
module ComputeNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_9] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h4;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_10] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: shl] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_11] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_12] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [63:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [63:0] io_idx_0_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] base_addr_R_data; // @[GepNode.scala 884:28]
  reg  base_addr_valid_R; // @[GepNode.scala 885:34]
  reg [63:0] idx_R_0_data; // @[GepNode.scala 888:39]
  reg  idx_valid_R_0; // @[GepNode.scala 889:45]
  reg  state; // @[GepNode.scala 893:22]
  wire  _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_11 | base_addr_valid_R; // @[GepNode.scala 909:31]
  wire  _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_13 | idx_valid_R_0; // @[GepNode.scala 916:28]
  wire [67:0] seek_value = idx_R_0_data * 64'h8; // @[GepNode.scala 924:21]
  wire [67:0] _GEN_52 = {{4'd0}, base_addr_R_data}; // @[GepNode.scala 932:35]
  wire [67:0] data_out = _GEN_52 + seek_value; // @[GepNode.scala 932:35]
  wire  _T_15 = ~state; // @[Conditional.scala 37:30]
  wire  _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 948:27]
  wire  _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 948:48]
  wire  _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _GEN_17 = _T_17 | state; // @[GepNode.scala 948:78]
  wire  _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_26 = ~reset; // @[GepNode.scala 968:17]
  wire  _GEN_53 = ~_T_15; // @[GepNode.scala 968:17]
  wire  _GEN_54 = _GEN_53 & state; // @[GepNode.scala 968:17]
  wire  _GEN_55 = _GEN_54 & _T_22; // @[GepNode.scala 968:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 194:21]
  assign io_Out_0_bits_data = data_out[63:0]; // @[GepNode.scala 936:25]
  assign io_baseAddress_ready = ~base_addr_valid_R; // @[GepNode.scala 908:24]
  assign io_idx_0_ready = ~idx_valid_R_0; // @[GepNode.scala 915:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  base_addr_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  idx_R_0_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_15) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_22) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_15) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_22) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      if (_T_17) begin
        out_valid_R_0 <= _T_19;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      base_addr_R_data <= 64'h0;
    end else if (_T_15) begin
      if (_T_11) begin
        base_addr_R_data <= io_baseAddress_bits_data;
      end
    end else if (state) begin
      if (_T_22) begin
        base_addr_R_data <= 64'h0;
      end else if (_T_11) begin
        base_addr_R_data <= io_baseAddress_bits_data;
      end
    end else if (_T_11) begin
      base_addr_R_data <= io_baseAddress_bits_data;
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else if (_T_15) begin
      base_addr_valid_R <= _GEN_11;
    end else if (state) begin
      if (_T_22) begin
        base_addr_valid_R <= 1'h0;
      end else begin
        base_addr_valid_R <= _GEN_11;
      end
    end else begin
      base_addr_valid_R <= _GEN_11;
    end
    if (reset) begin
      idx_R_0_data <= 64'h0;
    end else if (_T_15) begin
      if (_T_13) begin
        idx_R_0_data <= io_idx_0_bits_data;
      end
    end else if (state) begin
      if (_T_22) begin
        idx_R_0_data <= 64'h0;
      end else if (_T_13) begin
        idx_R_0_data <= io_idx_0_bits_data;
      end
    end else if (_T_13) begin
      idx_R_0_data <= io_idx_0_bits_data;
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      idx_valid_R_0 <= _GEN_15;
    end else if (state) begin
      if (_T_22) begin
        idx_valid_R_0 <= 1'h0;
      end else begin
        idx_valid_R_0 <= _GEN_15;
      end
    end else begin
      idx_valid_R_0 <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_15) begin
      state <= _GEN_17;
    end else if (state) begin
      if (_T_22) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [GEP] [Gep_arrayidx13] [Pred: %d][Out: 0x%x] [Cycle: %d]\n",enable_R_taskID,enable_R_control,data_out,cycleCount); // @[GepNode.scala 968:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoadCache(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [63:0] io_GepAddr_bits_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [63:0] io_MemReq_bits_addr,
  input         io_MemResp_valid,
  input  [63:0] io_MemResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_4 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 632:29]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [63:0] addr_R_data; // @[LoadCache.scala 58:23]
  reg  addr_valid_R; // @[LoadCache.scala 59:29]
  reg [63:0] data_R_data; // @[LoadCache.scala 62:23]
  reg [1:0] state; // @[LoadCache.scala 67:22]
  wire  _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | addr_valid_R; // @[LoadCache.scala 76:27]
  wire  _T_15 = enable_valid_R & addr_valid_R; // @[LoadCache.scala 95:20]
  wire  _T_16 = _T_15 & enable_R_control; // @[LoadCache.scala 95:36]
  wire  _T_23 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_24 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_25 = _T_23 | _T_24; // @[HandShaking.scala 725:29]
  wire  _T_44 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_49 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_25 = io_MemResp_valid | _GEN_1; // @[LoadCache.scala 214:30]
  wire  _T_51 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [14:0] _T_62 = value + 15'h1; // @[Counter.scala 39:22]
  wire  _T_64 = ~reset; // @[LoadCache.scala 254:17]
  wire  _GEN_78 = ~_T_44; // @[LoadCache.scala 254:17]
  wire  _GEN_79 = ~_T_50; // @[LoadCache.scala 254:17]
  wire  _GEN_80 = _GEN_78 & _GEN_79; // @[LoadCache.scala 254:17]
  wire  _GEN_81 = _GEN_80 & _T_51; // @[LoadCache.scala 254:17]
  wire  _GEN_82 = _GEN_81 & _T_25; // @[LoadCache.scala 254:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 630:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadCache.scala 158:20]
  assign io_GepAddr_ready = ~addr_valid_R; // @[LoadCache.scala 75:20]
  assign io_MemReq_valid = _T_44 & _T_16; // @[LoadCache.scala 162:19 LoadCache.scala 185:27]
  assign io_MemReq_bits_addr = addr_R_data; // @[LoadCache.scala 164:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[14:0];
  _RAND_7 = {2{`RANDOM}};
  addr_R_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  data_R_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_44) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_50) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_44) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_50) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_44) begin
      if (_T_15) begin
        if (enable_R_control) begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end else begin
          out_valid_R_0 <= _T_49;
        end
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_50) begin
      out_valid_R_0 <= _GEN_25;
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      value <= 15'h0;
    end else if (!(_T_44)) begin
      if (!(_T_50)) begin
        if (_T_51) begin
          if (_T_25) begin
            value <= _T_62;
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 64'h0;
    end else if (_T_44) begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_50) begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        addr_R_data <= 64'h0;
      end else if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_14) begin
      addr_R_data <= io_GepAddr_bits_data;
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else if (_T_44) begin
      addr_valid_R <= _GEN_11;
    end else if (_T_50) begin
      addr_valid_R <= _GEN_11;
    end else if (_T_51) begin
      if (_T_25) begin
        addr_valid_R <= 1'h0;
      end else begin
        addr_valid_R <= _GEN_11;
      end
    end else begin
      addr_valid_R <= _GEN_11;
    end
    if (reset) begin
      data_R_data <= 64'h0;
    end else if (!(_T_44)) begin
      if (_T_50) begin
        if (io_MemResp_valid) begin
          data_R_data <= io_MemResp_bits_data;
        end
      end else if (_T_51) begin
        if (_T_25) begin
          data_R_data <= 64'h0;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_44) begin
      if (_T_15) begin
        if (enable_R_control) begin
          if (io_MemReq_ready) begin
            state <= 2'h1;
          end
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_50) begin
      if (io_MemResp_valid) begin
        state <= 2'h2;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOAD] [ld_14] [Pred: %d] [Iter: %d] [Addr: %d] [Data: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,value,addr_R_data,data_R_data,cycleCount); // @[LoadCache.scala 254:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_4(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  state; // @[BranchNode.scala 588:22]
  wire  _T_11 = ~state; // @[Conditional.scala 37:30]
  wire  _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_16 = ~reset; // @[BranchNode.scala 616:17]
  wire  _GEN_8 = enable_valid_R | state; // @[BranchNode.scala 611:46]
  wire  _GEN_10 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 611:46]
  wire  _T_18 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_19 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_20 = _T_18 | _T_19; // @[HandShaking.scala 725:29]
  wire  _GEN_31 = _T_11 & enable_valid_R; // @[BranchNode.scala 616:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = _T_11 ? _GEN_10 : out_valid_R_0; // @[HandShaking.scala 630:21 BranchNode.scala 614:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 607:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 607:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_R_control <= 1'h0;
      end else if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_11) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_20) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_20) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_11) begin
      if (enable_valid_R) begin
        out_valid_R_0 <= _T_14;
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_11) begin
      state <= _GEN_8;
    end else if (state) begin
      if (_T_20) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_31 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [UBR] [br_15] [Out: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,cycleCount); // @[BranchNode.scala 616:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [63:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [63:0] io_Out_2_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] in_data_R_1_data; // @[PhiNode.scala 203:26]
  reg  in_data_valid_R_0; // @[PhiNode.scala 204:32]
  reg  in_data_valid_R_1; // @[PhiNode.scala 204:32]
  reg  enable_R_control; // @[PhiNode.scala 207:25]
  reg  enable_valid_R; // @[PhiNode.scala 208:31]
  reg [1:0] mask_R; // @[PhiNode.scala 211:23]
  reg  mask_valid_R; // @[PhiNode.scala 212:29]
  reg [1:0] state; // @[PhiNode.scala 216:22]
  reg  out_valid_R_0; // @[PhiNode.scala 219:49]
  reg  out_valid_R_1; // @[PhiNode.scala 219:49]
  reg  out_valid_R_2; // @[PhiNode.scala 219:49]
  reg  fire_R_0; // @[PhiNode.scala 221:44]
  reg  fire_R_1; // @[PhiNode.scala 221:44]
  reg  fire_R_2; // @[PhiNode.scala 221:44]
  wire  _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_3 = _T_10 | mask_valid_R; // @[PhiNode.scala 239:24]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_7 = _T_12 | enable_valid_R; // @[PhiNode.scala 246:26]
  wire  _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 254:29]
  wire  _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 254:29]
  wire [1:0] _T_19 = {mask_R[0],mask_R[1]}; // @[Cat.scala 29:58]
  wire  sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  wire  _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_16 = _T_20 | fire_R_0; // @[PhiNode.scala 276:26]
  wire  _GEN_17 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 276:26]
  wire  _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = _T_21 | fire_R_1; // @[PhiNode.scala 276:26]
  wire  _GEN_19 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 276:26]
  wire  _T_22 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_20 = _T_22 | fire_R_2; // @[PhiNode.scala 276:26]
  wire  _GEN_21 = _T_22 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 276:26]
  wire  fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 283:74]
  wire  fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 283:74]
  wire  fire_mask_2 = fire_R_2 | _T_22; // @[PhiNode.scala 283:74]
  wire [63:0] _GEN_28 = sel ? in_data_R_1_data : 64'h0; // @[PhiNode.scala 312:12]
  wire  _T_31 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 286:30]
  wire  _T_32 = enable_valid_R & _T_31; // @[PhiNode.scala 290:20]
  wire  _T_37 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_42 = ~reset; // @[PhiNode.scala 350:19]
  wire [4:0] _GEN_37 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 350:19]
  wire  _GEN_40 = _T_32 | _GEN_17; // @[PhiNode.scala 327:66]
  wire  _GEN_41 = _T_32 | _GEN_19; // @[PhiNode.scala 327:66]
  wire  _GEN_42 = _T_32 | _GEN_21; // @[PhiNode.scala 327:66]
  wire  _T_45 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_46 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 364:31]
  wire  _T_47 = _T_46 & fire_mask_2; // @[PhiNode.scala 364:31]
  wire  _T_51 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_81 = _T_51 ? 64'h0 : _GEN_28; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_127 = _T_45 ? _GEN_28 : _GEN_81; // @[Conditional.scala 39:67]
  wire  _GEN_167 = _T_37 & _T_32; // @[PhiNode.scala 350:19]
  wire  _GEN_168 = _GEN_167 & enable_R_control; // @[PhiNode.scala 350:19]
  wire  _GEN_170 = ~enable_R_control; // @[PhiNode.scala 357:19]
  wire  _GEN_171 = _GEN_167 & _GEN_170; // @[PhiNode.scala 357:19]
  assign io_enable_ready = ~enable_valid_R; // @[PhiNode.scala 245:19]
  assign io_InData_0_ready = ~in_data_valid_R_0; // @[PhiNode.scala 253:24]
  assign io_InData_1_ready = ~in_data_valid_R_1; // @[PhiNode.scala 253:24]
  assign io_Mask_ready = ~mask_valid_R; // @[PhiNode.scala 238:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 322:21]
  assign io_Out_0_bits_data = _T_37 ? _GEN_28 : _GEN_127; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 322:21]
  assign io_Out_1_bits_data = _T_37 ? _GEN_28 : _GEN_127; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 322:21]
  assign io_Out_2_bits_data = _T_37 ? _GEN_28 : _GEN_127; // @[PhiNode.scala 321:20 PhiNode.scala 392:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {2{`RANDOM}};
  in_data_R_1_data = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_R_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fire_R_2 = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      in_data_R_1_data <= 64'h0;
    end else if (_T_37) begin
      if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_45) begin
      if (_T_47) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        in_data_R_1_data <= 64'h0;
      end else if (_T_16) begin
        in_data_R_1_data <= io_InData_1_bits_data;
      end
    end else if (_T_16) begin
      in_data_R_1_data <= io_InData_1_bits_data;
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      in_data_valid_R_0 <= _GEN_11;
    end else if (_T_45) begin
      if (_T_47) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        in_data_valid_R_0 <= 1'h0;
      end else begin
        in_data_valid_R_0 <= _GEN_11;
      end
    end else begin
      in_data_valid_R_0 <= _GEN_11;
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else if (_T_37) begin
      in_data_valid_R_1 <= _GEN_15;
    end else if (_T_45) begin
      if (_T_47) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        in_data_valid_R_1 <= 1'h0;
      end else begin
        in_data_valid_R_1 <= _GEN_15;
      end
    end else begin
      in_data_valid_R_1 <= _GEN_15;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_37) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_45) begin
      if (_T_47) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_37) begin
      enable_valid_R <= _GEN_7;
    end else if (_T_45) begin
      if (_T_47) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_7;
      end
    end else begin
      enable_valid_R <= _GEN_7;
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else if (_T_37) begin
      if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_45) begin
      if (_T_47) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        mask_R <= 2'h0;
      end else if (_T_10) begin
        mask_R <= io_Mask_bits;
      end
    end else if (_T_10) begin
      mask_R <= io_Mask_bits;
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else if (_T_37) begin
      mask_valid_R <= _GEN_3;
    end else if (_T_45) begin
      if (_T_47) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        mask_valid_R <= 1'h0;
      end else begin
        mask_valid_R <= _GEN_3;
      end
    end else begin
      mask_valid_R <= _GEN_3;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_37) begin
      if (_T_32) begin
        if (enable_R_control) begin
          state <= 2'h1;
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_45) begin
      if (_T_47) begin
        state <= 2'h0;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        state <= 2'h0;
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_0 <= _GEN_40;
    end else if (_T_20) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_1 <= _GEN_41;
    end else if (_T_21) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else if (_T_37) begin
      out_valid_R_2 <= _GEN_42;
    end else if (_T_22) begin
      out_valid_R_2 <= 1'h0;
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else if (_T_37) begin
      fire_R_0 <= _GEN_16;
    end else if (_T_45) begin
      if (_T_47) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        fire_R_0 <= 1'h0;
      end else begin
        fire_R_0 <= _GEN_16;
      end
    end else begin
      fire_R_0 <= _GEN_16;
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else if (_T_37) begin
      fire_R_1 <= _GEN_18;
    end else if (_T_45) begin
      if (_T_47) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        fire_R_1 <= 1'h0;
      end else begin
        fire_R_1 <= _GEN_18;
      end
    end else begin
      fire_R_1 <= _GEN_18;
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else if (_T_37) begin
      fire_R_2 <= _GEN_20;
    end else if (_T_45) begin
      if (_T_47) begin
        fire_R_2 <= 1'h0;
      end else begin
        fire_R_2 <= _GEN_20;
      end
    end else if (_T_51) begin
      if (_T_47) begin
        fire_R_2 <= 1'h0;
      end else begin
        fire_R_2 <= _GEN_20;
      end
    end else begin
      fire_R_2 <= _GEN_20;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_168 & _T_42) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv16] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_37,enable_R_control,_GEN_28,cycleCount); // @[PhiNode.scala 350:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_171 & _T_42) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [PHI] [phiindvars_iv16] [Pred: %d] [Out: %d] [Cycle: %d]\n",_GEN_37,enable_R_control,_GEN_28,cycleCount); // @[PhiNode.scala 357:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_17] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_18] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [63:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [63:0] io_idx_0_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] base_addr_R_data; // @[GepNode.scala 884:28]
  reg  base_addr_valid_R; // @[GepNode.scala 885:34]
  reg [63:0] idx_R_0_data; // @[GepNode.scala 888:39]
  reg  idx_valid_R_0; // @[GepNode.scala 889:45]
  reg  state; // @[GepNode.scala 893:22]
  wire  _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_11 | base_addr_valid_R; // @[GepNode.scala 909:31]
  wire  _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_13 | idx_valid_R_0; // @[GepNode.scala 916:28]
  wire [67:0] seek_value = idx_R_0_data * 64'h8; // @[GepNode.scala 924:21]
  wire [67:0] _GEN_52 = {{4'd0}, base_addr_R_data}; // @[GepNode.scala 932:35]
  wire [67:0] data_out = _GEN_52 + seek_value; // @[GepNode.scala 932:35]
  wire  _T_15 = ~state; // @[Conditional.scala 37:30]
  wire  _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 948:27]
  wire  _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 948:48]
  wire  _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _GEN_17 = _T_17 | state; // @[GepNode.scala 948:78]
  wire  _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_26 = ~reset; // @[GepNode.scala 968:17]
  wire  _GEN_53 = ~_T_15; // @[GepNode.scala 968:17]
  wire  _GEN_54 = _GEN_53 & state; // @[GepNode.scala 968:17]
  wire  _GEN_55 = _GEN_54 & _T_22; // @[GepNode.scala 968:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 194:21]
  assign io_Out_0_bits_data = data_out[63:0]; // @[GepNode.scala 936:25]
  assign io_baseAddress_ready = ~base_addr_valid_R; // @[GepNode.scala 908:24]
  assign io_idx_0_ready = ~idx_valid_R_0; // @[GepNode.scala 915:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  base_addr_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  idx_R_0_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_15) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_22) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_15) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_22) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      if (_T_17) begin
        out_valid_R_0 <= _T_19;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      base_addr_R_data <= 64'h0;
    end else if (_T_15) begin
      if (_T_11) begin
        base_addr_R_data <= io_baseAddress_bits_data;
      end
    end else if (state) begin
      if (_T_22) begin
        base_addr_R_data <= 64'h0;
      end else if (_T_11) begin
        base_addr_R_data <= io_baseAddress_bits_data;
      end
    end else if (_T_11) begin
      base_addr_R_data <= io_baseAddress_bits_data;
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else if (_T_15) begin
      base_addr_valid_R <= _GEN_11;
    end else if (state) begin
      if (_T_22) begin
        base_addr_valid_R <= 1'h0;
      end else begin
        base_addr_valid_R <= _GEN_11;
      end
    end else begin
      base_addr_valid_R <= _GEN_11;
    end
    if (reset) begin
      idx_R_0_data <= 64'h0;
    end else if (_T_15) begin
      if (_T_13) begin
        idx_R_0_data <= io_idx_0_bits_data;
      end
    end else if (state) begin
      if (_T_22) begin
        idx_R_0_data <= 64'h0;
      end else if (_T_13) begin
        idx_R_0_data <= io_idx_0_bits_data;
      end
    end else if (_T_13) begin
      idx_R_0_data <= io_idx_0_bits_data;
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else if (_T_15) begin
      idx_valid_R_0 <= _GEN_15;
    end else if (state) begin
      if (_T_22) begin
        idx_valid_R_0 <= 1'h0;
      end else begin
        idx_valid_R_0 <= _GEN_15;
      end
    end else begin
      idx_valid_R_0 <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_15) begin
      state <= _GEN_17;
    end else if (state) begin
      if (_T_22) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [GEP] [Gep_arrayidx2019] [Pred: %d][Out: 0x%x] [Cycle: %d]\n",enable_R_taskID,enable_R_control,data_out,cycleCount); // @[GepNode.scala 968:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoadCache_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [63:0] io_GepAddr_bits_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [63:0] io_MemReq_bits_addr,
  input         io_MemResp_valid,
  input  [63:0] io_MemResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_4 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 632:29]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [63:0] addr_R_data; // @[LoadCache.scala 58:23]
  reg  addr_valid_R; // @[LoadCache.scala 59:29]
  reg [63:0] data_R_data; // @[LoadCache.scala 62:23]
  reg [1:0] state; // @[LoadCache.scala 67:22]
  wire  _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | addr_valid_R; // @[LoadCache.scala 76:27]
  wire  _T_15 = enable_valid_R & addr_valid_R; // @[LoadCache.scala 95:20]
  wire  _T_16 = _T_15 & enable_R_control; // @[LoadCache.scala 95:36]
  wire  _T_23 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_24 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_25 = _T_23 | _T_24; // @[HandShaking.scala 725:29]
  wire  _T_44 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_49 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_25 = io_MemResp_valid | _GEN_1; // @[LoadCache.scala 214:30]
  wire  _T_51 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [14:0] _T_62 = value + 15'h1; // @[Counter.scala 39:22]
  wire  _T_64 = ~reset; // @[LoadCache.scala 254:17]
  wire  _GEN_78 = ~_T_44; // @[LoadCache.scala 254:17]
  wire  _GEN_79 = ~_T_50; // @[LoadCache.scala 254:17]
  wire  _GEN_80 = _GEN_78 & _GEN_79; // @[LoadCache.scala 254:17]
  wire  _GEN_81 = _GEN_80 & _T_51; // @[LoadCache.scala 254:17]
  wire  _GEN_82 = _GEN_81 & _T_25; // @[LoadCache.scala 254:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 630:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadCache.scala 158:20]
  assign io_GepAddr_ready = ~addr_valid_R; // @[LoadCache.scala 75:20]
  assign io_MemReq_valid = _T_44 & _T_16; // @[LoadCache.scala 162:19 LoadCache.scala 185:27]
  assign io_MemReq_bits_addr = addr_R_data; // @[LoadCache.scala 164:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[14:0];
  _RAND_7 = {2{`RANDOM}};
  addr_R_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  data_R_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_44) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_50) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_44) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_50) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_44) begin
      if (_T_15) begin
        if (enable_R_control) begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end else begin
          out_valid_R_0 <= _T_49;
        end
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_50) begin
      out_valid_R_0 <= _GEN_25;
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      value <= 15'h0;
    end else if (!(_T_44)) begin
      if (!(_T_50)) begin
        if (_T_51) begin
          if (_T_25) begin
            value <= _T_62;
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 64'h0;
    end else if (_T_44) begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_50) begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        addr_R_data <= 64'h0;
      end else if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_14) begin
      addr_R_data <= io_GepAddr_bits_data;
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else if (_T_44) begin
      addr_valid_R <= _GEN_11;
    end else if (_T_50) begin
      addr_valid_R <= _GEN_11;
    end else if (_T_51) begin
      if (_T_25) begin
        addr_valid_R <= 1'h0;
      end else begin
        addr_valid_R <= _GEN_11;
      end
    end else begin
      addr_valid_R <= _GEN_11;
    end
    if (reset) begin
      data_R_data <= 64'h0;
    end else if (!(_T_44)) begin
      if (_T_50) begin
        if (io_MemResp_valid) begin
          data_R_data <= io_MemResp_bits_data;
        end
      end else if (_T_51) begin
        if (_T_25) begin
          data_R_data <= 64'h0;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_44) begin
      if (_T_15) begin
        if (enable_R_control) begin
          if (io_MemReq_ready) begin
            state <= 2'h1;
          end
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_50) begin
      if (io_MemResp_valid) begin
        state <= 2'h2;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOAD] [ld_20] [Pred: %d] [Iter: %d] [Addr: %d] [Data: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,value,addr_R_data,data_R_data,cycleCount); // @[LoadCache.scala 254:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module RoundAnyRawFNToRecFN(
  input         io_in_isZero,
  input  [8:0]  io_in_sExp,
  input  [64:0] io_in_sig,
  output [64:0] io_out
);
  wire [11:0] _GEN_0 = {{3{io_in_sExp[8]}},io_in_sExp}; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] _T_3 = $signed(_GEN_0) + 12'sh780; // @[RoundAnyRawFNToRecFN.scala 102:25]
  wire [12:0] sAdjustedExp = {1'b0,$signed(_T_3[11:0])}; // @[RoundAnyRawFNToRecFN.scala 104:31]
  wire  _T_7 = |io_in_sig[9:0]; // @[RoundAnyRawFNToRecFN.scala 115:60]
  wire [55:0] adjustedSig = {io_in_sig[64:10],_T_7}; // @[Cat.scala 29:58]
  wire [55:0] _T_14 = adjustedSig & 56'h2; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_15 = |_T_14; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_16 = adjustedSig & 56'h1; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_17 = |_T_16; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  common_inexact = _T_15 | _T_17; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire [55:0] _T_34 = adjustedSig & 56'hfffffffffffffc; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [54:0] _T_38 = common_inexact ? 55'h1 : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_1 = {{1'd0}, _T_34[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_39 = _GEN_1 | _T_38; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [2:0] _T_42 = {1'b0,$signed(_T_39[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_2 = {{10{_T_42[2]}},_T_42}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_43 = $signed(sAdjustedExp) + $signed(_GEN_2); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut = _T_43[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut = _T_39[51:0]; // @[RoundAnyRawFNToRecFN.scala 189:27]
  wire [11:0] _T_75 = io_in_isZero ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _T_76 = ~_T_75; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [11:0] expOut = common_expOut & _T_76; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [51:0] fractOut = io_in_isZero ? 52'h0 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [12:0] _T_101 = {1'h0,expOut}; // @[Cat.scala 29:58]
  assign io_out = {_T_101,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
endmodule
module INToRecFN(
  input  [63:0] io_in,
  output [64:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[INToRecFN.scala 59:15]
  wire [8:0] roundAnyRawFNToRecFN_io_in_sExp; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_in_sig; // @[INToRecFN.scala 59:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 59:15]
  wire [127:0] _T_5 = {64'h0,io_in}; // @[Cat.scala 29:58]
  wire [5:0] _T_71 = _T_5[1] ? 6'h3e : 6'h3f; // @[Mux.scala 47:69]
  wire [5:0] _T_72 = _T_5[2] ? 6'h3d : _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_73 = _T_5[3] ? 6'h3c : _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_74 = _T_5[4] ? 6'h3b : _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_75 = _T_5[5] ? 6'h3a : _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_76 = _T_5[6] ? 6'h39 : _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_77 = _T_5[7] ? 6'h38 : _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_78 = _T_5[8] ? 6'h37 : _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_79 = _T_5[9] ? 6'h36 : _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_80 = _T_5[10] ? 6'h35 : _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_81 = _T_5[11] ? 6'h34 : _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_82 = _T_5[12] ? 6'h33 : _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_83 = _T_5[13] ? 6'h32 : _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_84 = _T_5[14] ? 6'h31 : _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_85 = _T_5[15] ? 6'h30 : _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_86 = _T_5[16] ? 6'h2f : _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_87 = _T_5[17] ? 6'h2e : _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_88 = _T_5[18] ? 6'h2d : _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_89 = _T_5[19] ? 6'h2c : _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_90 = _T_5[20] ? 6'h2b : _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_91 = _T_5[21] ? 6'h2a : _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_92 = _T_5[22] ? 6'h29 : _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_93 = _T_5[23] ? 6'h28 : _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_94 = _T_5[24] ? 6'h27 : _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_95 = _T_5[25] ? 6'h26 : _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_96 = _T_5[26] ? 6'h25 : _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_97 = _T_5[27] ? 6'h24 : _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_98 = _T_5[28] ? 6'h23 : _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_99 = _T_5[29] ? 6'h22 : _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_100 = _T_5[30] ? 6'h21 : _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_101 = _T_5[31] ? 6'h20 : _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_102 = _T_5[32] ? 6'h1f : _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_103 = _T_5[33] ? 6'h1e : _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_104 = _T_5[34] ? 6'h1d : _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_105 = _T_5[35] ? 6'h1c : _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_106 = _T_5[36] ? 6'h1b : _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_107 = _T_5[37] ? 6'h1a : _T_106; // @[Mux.scala 47:69]
  wire [5:0] _T_108 = _T_5[38] ? 6'h19 : _T_107; // @[Mux.scala 47:69]
  wire [5:0] _T_109 = _T_5[39] ? 6'h18 : _T_108; // @[Mux.scala 47:69]
  wire [5:0] _T_110 = _T_5[40] ? 6'h17 : _T_109; // @[Mux.scala 47:69]
  wire [5:0] _T_111 = _T_5[41] ? 6'h16 : _T_110; // @[Mux.scala 47:69]
  wire [5:0] _T_112 = _T_5[42] ? 6'h15 : _T_111; // @[Mux.scala 47:69]
  wire [5:0] _T_113 = _T_5[43] ? 6'h14 : _T_112; // @[Mux.scala 47:69]
  wire [5:0] _T_114 = _T_5[44] ? 6'h13 : _T_113; // @[Mux.scala 47:69]
  wire [5:0] _T_115 = _T_5[45] ? 6'h12 : _T_114; // @[Mux.scala 47:69]
  wire [5:0] _T_116 = _T_5[46] ? 6'h11 : _T_115; // @[Mux.scala 47:69]
  wire [5:0] _T_117 = _T_5[47] ? 6'h10 : _T_116; // @[Mux.scala 47:69]
  wire [5:0] _T_118 = _T_5[48] ? 6'hf : _T_117; // @[Mux.scala 47:69]
  wire [5:0] _T_119 = _T_5[49] ? 6'he : _T_118; // @[Mux.scala 47:69]
  wire [5:0] _T_120 = _T_5[50] ? 6'hd : _T_119; // @[Mux.scala 47:69]
  wire [5:0] _T_121 = _T_5[51] ? 6'hc : _T_120; // @[Mux.scala 47:69]
  wire [5:0] _T_122 = _T_5[52] ? 6'hb : _T_121; // @[Mux.scala 47:69]
  wire [5:0] _T_123 = _T_5[53] ? 6'ha : _T_122; // @[Mux.scala 47:69]
  wire [5:0] _T_124 = _T_5[54] ? 6'h9 : _T_123; // @[Mux.scala 47:69]
  wire [5:0] _T_125 = _T_5[55] ? 6'h8 : _T_124; // @[Mux.scala 47:69]
  wire [5:0] _T_126 = _T_5[56] ? 6'h7 : _T_125; // @[Mux.scala 47:69]
  wire [5:0] _T_127 = _T_5[57] ? 6'h6 : _T_126; // @[Mux.scala 47:69]
  wire [5:0] _T_128 = _T_5[58] ? 6'h5 : _T_127; // @[Mux.scala 47:69]
  wire [5:0] _T_129 = _T_5[59] ? 6'h4 : _T_128; // @[Mux.scala 47:69]
  wire [5:0] _T_130 = _T_5[60] ? 6'h3 : _T_129; // @[Mux.scala 47:69]
  wire [5:0] _T_131 = _T_5[61] ? 6'h2 : _T_130; // @[Mux.scala 47:69]
  wire [5:0] _T_132 = _T_5[62] ? 6'h1 : _T_131; // @[Mux.scala 47:69]
  wire [5:0] _T_133 = _T_5[63] ? 6'h0 : _T_132; // @[Mux.scala 47:69]
  wire [126:0] _GEN_0 = {{63'd0}, _T_5[63:0]}; // @[rawFloatFromIN.scala 55:22]
  wire [126:0] _T_134 = _GEN_0 << _T_133; // @[rawFloatFromIN.scala 55:22]
  wire [5:0] _T_139 = ~_T_133; // @[rawFloatFromIN.scala 63:39]
  wire [7:0] _T_140 = {2'h2,_T_139}; // @[Cat.scala 29:58]
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN ( // @[INToRecFN.scala 59:15]
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[INToRecFN.scala 72:23]
  assign roundAnyRawFNToRecFN_io_in_isZero = ~_T_134[63]; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = {1'b0,$signed(_T_140)}; // @[INToRecFN.scala 69:44]
  assign roundAnyRawFNToRecFN_io_in_sig = {{1'd0}, _T_134[63:0]}; // @[INToRecFN.scala 69:44]
endmodule
module MulAddRecFNToRaw_preMul(
  input  [64:0]  io_a,
  input  [64:0]  io_b,
  input  [64:0]  io_c,
  output [52:0]  io_mulAddA,
  output [52:0]  io_mulAddB,
  output [105:0] io_mulAddC,
  output         io_toPostMul_isSigNaNAny,
  output         io_toPostMul_isNaNAOrB,
  output         io_toPostMul_isInfA,
  output         io_toPostMul_isZeroA,
  output         io_toPostMul_isInfB,
  output         io_toPostMul_isZeroB,
  output         io_toPostMul_signProd,
  output         io_toPostMul_isNaNC,
  output         io_toPostMul_isInfC,
  output         io_toPostMul_isZeroC,
  output [12:0]  io_toPostMul_sExpSum,
  output         io_toPostMul_doSubMags,
  output         io_toPostMul_CIsDominant,
  output [5:0]   io_toPostMul_CDom_CAlignDist,
  output [54:0]  io_toPostMul_highAlignedSigC,
  output         io_toPostMul_bit0AlignedSigC
);
  wire  rawA_isZero = io_a[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_4 = io_a[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawA_isNaN = _T_4 & io_a[61]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_8 = ~io_a[61]; // @[rawFloatFromRecFN.scala 56:36]
  wire  rawA_sign = io_a[64]; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawA_sExp = {1'b0,$signed(io_a[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _T_12 = ~rawA_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [53:0] rawA_sig = {1'h0,_T_12,io_a[51:0]}; // @[Cat.scala 29:58]
  wire  rawB_isZero = io_b[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_20 = io_b[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawB_isNaN = _T_20 & io_b[61]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_24 = ~io_b[61]; // @[rawFloatFromRecFN.scala 56:36]
  wire  rawB_sign = io_b[64]; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawB_sExp = {1'b0,$signed(io_b[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _T_28 = ~rawB_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [53:0] rawB_sig = {1'h0,_T_28,io_b[51:0]}; // @[Cat.scala 29:58]
  wire  rawC_isZero = io_c[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_36 = io_c[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  rawC_isNaN = _T_36 & io_c[61]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_40 = ~io_c[61]; // @[rawFloatFromRecFN.scala 56:36]
  wire  rawC_sign = io_c[64]; // @[rawFloatFromRecFN.scala 58:25]
  wire [12:0] rawC_sExp = {1'b0,$signed(io_c[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _T_44 = ~rawC_isZero; // @[rawFloatFromRecFN.scala 60:39]
  wire [53:0] rawC_sig = {1'h0,_T_44,io_c[51:0]}; // @[Cat.scala 29:58]
  wire  signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 98:30]
  wire [13:0] _T_50 = $signed(rawA_sExp) + $signed(rawB_sExp); // @[MulAddRecFN.scala 101:19]
  wire [13:0] sExpAlignedProd = $signed(_T_50) - 14'sh7c8; // @[MulAddRecFN.scala 101:32]
  wire  doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 103:30]
  wire [13:0] _GEN_0 = {{1{rawC_sExp[12]}},rawC_sExp}; // @[MulAddRecFN.scala 107:42]
  wire [13:0] sNatCAlignDist = $signed(sExpAlignedProd) - $signed(_GEN_0); // @[MulAddRecFN.scala 107:42]
  wire [12:0] posNatCAlignDist = sNatCAlignDist[12:0]; // @[MulAddRecFN.scala 108:42]
  wire  _T_57 = rawA_isZero | rawB_isZero; // @[MulAddRecFN.scala 109:35]
  wire  _T_58 = $signed(sNatCAlignDist) < 14'sh0; // @[MulAddRecFN.scala 109:69]
  wire  isMinCAlign = _T_57 | _T_58; // @[MulAddRecFN.scala 109:50]
  wire  _T_60 = posNatCAlignDist <= 13'h35; // @[MulAddRecFN.scala 111:60]
  wire  _T_61 = isMinCAlign | _T_60; // @[MulAddRecFN.scala 111:39]
  wire  CIsDominant = _T_44 & _T_61; // @[MulAddRecFN.scala 111:23]
  wire  _T_62 = posNatCAlignDist < 13'ha1; // @[MulAddRecFN.scala 115:34]
  wire [7:0] _T_64 = _T_62 ? posNatCAlignDist[7:0] : 8'ha1; // @[MulAddRecFN.scala 115:16]
  wire [7:0] CAlignDist = isMinCAlign ? 8'h0 : _T_64; // @[MulAddRecFN.scala 113:12]
  wire [53:0] _T_65 = ~rawC_sig; // @[MulAddRecFN.scala 121:28]
  wire [53:0] _T_66 = doSubMags ? _T_65 : rawC_sig; // @[MulAddRecFN.scala 121:16]
  wire [110:0] _T_68 = doSubMags ? 111'h7fffffffffffffffffffffffffff : 111'h0; // @[Bitwise.scala 72:12]
  wire [164:0] _T_70 = {_T_66,_T_68}; // @[MulAddRecFN.scala 123:11]
  wire [164:0] mainAlignedSigC = $signed(_T_70) >>> CAlignDist; // @[MulAddRecFN.scala 123:17]
  wire  _T_74 = |rawC_sig[3:0]; // @[primitives.scala 121:54]
  wire  _T_76 = |rawC_sig[7:4]; // @[primitives.scala 121:54]
  wire  _T_78 = |rawC_sig[11:8]; // @[primitives.scala 121:54]
  wire  _T_80 = |rawC_sig[15:12]; // @[primitives.scala 121:54]
  wire  _T_82 = |rawC_sig[19:16]; // @[primitives.scala 121:54]
  wire  _T_84 = |rawC_sig[23:20]; // @[primitives.scala 121:54]
  wire  _T_86 = |rawC_sig[27:24]; // @[primitives.scala 121:54]
  wire  _T_88 = |rawC_sig[31:28]; // @[primitives.scala 121:54]
  wire  _T_90 = |rawC_sig[35:32]; // @[primitives.scala 121:54]
  wire  _T_92 = |rawC_sig[39:36]; // @[primitives.scala 121:54]
  wire  _T_94 = |rawC_sig[43:40]; // @[primitives.scala 121:54]
  wire  _T_96 = |rawC_sig[47:44]; // @[primitives.scala 121:54]
  wire  _T_98 = |rawC_sig[51:48]; // @[primitives.scala 121:54]
  wire  _T_100 = |rawC_sig[53:52]; // @[primitives.scala 124:57]
  wire [6:0] _T_106 = {_T_86,_T_84,_T_82,_T_80,_T_78,_T_76,_T_74}; // @[primitives.scala 125:20]
  wire [13:0] _T_113 = {_T_100,_T_98,_T_96,_T_94,_T_92,_T_90,_T_88,_T_106}; // @[primitives.scala 125:20]
  wire [64:0] _T_115 = -65'sh10000000000000000 >>> CAlignDist[7:2]; // @[primitives.scala 77:58]
  wire [7:0] _T_121 = {{4'd0}, _T_115[31:28]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_123 = {_T_115[27:24], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_125 = _T_123 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_126 = _T_121 | _T_125; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_1 = {{2'd0}, _T_126[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_131 = _GEN_1 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_133 = {_T_126[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_135 = _T_133 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_136 = _T_131 | _T_135; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2 = {{1'd0}, _T_136[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_141 = _GEN_2 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_143 = {_T_136[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_145 = _T_143 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_146 = _T_141 | _T_145; // @[Bitwise.scala 103:39]
  wire [12:0] _T_160 = {_T_146,_T_115[32],_T_115[33],_T_115[34],_T_115[35],_T_115[36]}; // @[Cat.scala 29:58]
  wire [13:0] _GEN_3 = {{1'd0}, _T_160}; // @[MulAddRecFN.scala 125:68]
  wire [13:0] _T_161 = _T_113 & _GEN_3; // @[MulAddRecFN.scala 125:68]
  wire  reduced4CExtra = |_T_161; // @[MulAddRecFN.scala 133:11]
  wire  _T_164 = &mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 137:39]
  wire  _T_165 = ~reduced4CExtra; // @[MulAddRecFN.scala 137:47]
  wire  _T_166 = _T_164 & _T_165; // @[MulAddRecFN.scala 137:44]
  wire  _T_168 = |mainAlignedSigC[2:0]; // @[MulAddRecFN.scala 138:39]
  wire  _T_169 = _T_168 | reduced4CExtra; // @[MulAddRecFN.scala 138:44]
  wire  _T_170 = doSubMags ? _T_166 : _T_169; // @[MulAddRecFN.scala 136:16]
  wire [161:0] _T_171 = mainAlignedSigC[164:3]; // @[Cat.scala 29:58]
  wire [162:0] alignedSigC = {_T_171,_T_170}; // @[Cat.scala 29:58]
  wire  _T_174 = ~rawA_sig[51]; // @[common.scala 81:49]
  wire  _T_175 = rawA_isNaN & _T_174; // @[common.scala 81:46]
  wire  _T_177 = ~rawB_sig[51]; // @[common.scala 81:49]
  wire  _T_178 = rawB_isNaN & _T_177; // @[common.scala 81:46]
  wire  _T_179 = _T_175 | _T_178; // @[MulAddRecFN.scala 149:32]
  wire  _T_181 = ~rawC_sig[51]; // @[common.scala 81:49]
  wire  _T_182 = rawC_isNaN & _T_181; // @[common.scala 81:46]
  wire [13:0] _T_187 = $signed(sExpAlignedProd) - 14'sh35; // @[MulAddRecFN.scala 161:53]
  wire [13:0] _T_188 = CIsDominant ? $signed({{1{rawC_sExp[12]}},rawC_sExp}) : $signed(_T_187); // @[MulAddRecFN.scala 161:12]
  assign io_mulAddA = rawA_sig[52:0]; // @[MulAddRecFN.scala 144:16]
  assign io_mulAddB = rawB_sig[52:0]; // @[MulAddRecFN.scala 145:16]
  assign io_mulAddC = alignedSigC[106:1]; // @[MulAddRecFN.scala 146:16]
  assign io_toPostMul_isSigNaNAny = _T_179 | _T_182; // @[MulAddRecFN.scala 148:30]
  assign io_toPostMul_isNaNAOrB = rawA_isNaN | rawB_isNaN; // @[MulAddRecFN.scala 151:28]
  assign io_toPostMul_isInfA = _T_4 & _T_8; // @[MulAddRecFN.scala 152:28]
  assign io_toPostMul_isZeroA = io_a[63:61] == 3'h0; // @[MulAddRecFN.scala 153:28]
  assign io_toPostMul_isInfB = _T_20 & _T_24; // @[MulAddRecFN.scala 154:28]
  assign io_toPostMul_isZeroB = io_b[63:61] == 3'h0; // @[MulAddRecFN.scala 155:28]
  assign io_toPostMul_signProd = rawA_sign ^ rawB_sign; // @[MulAddRecFN.scala 156:28]
  assign io_toPostMul_isNaNC = _T_36 & io_c[61]; // @[MulAddRecFN.scala 157:28]
  assign io_toPostMul_isInfC = _T_36 & _T_40; // @[MulAddRecFN.scala 158:28]
  assign io_toPostMul_isZeroC = io_c[63:61] == 3'h0; // @[MulAddRecFN.scala 159:28]
  assign io_toPostMul_sExpSum = _T_188[12:0]; // @[MulAddRecFN.scala 160:28]
  assign io_toPostMul_doSubMags = signProd ^ rawC_sign; // @[MulAddRecFN.scala 162:28]
  assign io_toPostMul_CIsDominant = _T_44 & _T_61; // @[MulAddRecFN.scala 163:30]
  assign io_toPostMul_CDom_CAlignDist = CAlignDist[5:0]; // @[MulAddRecFN.scala 164:34]
  assign io_toPostMul_highAlignedSigC = alignedSigC[161:107]; // @[MulAddRecFN.scala 165:34]
  assign io_toPostMul_bit0AlignedSigC = alignedSigC[0]; // @[MulAddRecFN.scala 167:34]
endmodule
module MulAddRecFNToRaw_postMul(
  input          io_fromPreMul_isSigNaNAny,
  input          io_fromPreMul_isNaNAOrB,
  input          io_fromPreMul_isInfA,
  input          io_fromPreMul_isZeroA,
  input          io_fromPreMul_isInfB,
  input          io_fromPreMul_isZeroB,
  input          io_fromPreMul_signProd,
  input          io_fromPreMul_isNaNC,
  input          io_fromPreMul_isInfC,
  input          io_fromPreMul_isZeroC,
  input  [12:0]  io_fromPreMul_sExpSum,
  input          io_fromPreMul_doSubMags,
  input          io_fromPreMul_CIsDominant,
  input  [5:0]   io_fromPreMul_CDom_CAlignDist,
  input  [54:0]  io_fromPreMul_highAlignedSigC,
  input          io_fromPreMul_bit0AlignedSigC,
  input  [106:0] io_mulAddResult,
  output         io_invalidExc,
  output         io_rawOut_isNaN,
  output         io_rawOut_isInf,
  output         io_rawOut_isZero,
  output         io_rawOut_sign,
  output [12:0]  io_rawOut_sExp,
  output [55:0]  io_rawOut_sig
);
  wire  CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 192:42]
  wire [54:0] _T_2 = io_fromPreMul_highAlignedSigC + 55'h1; // @[MulAddRecFN.scala 195:47]
  wire [54:0] _T_3 = io_mulAddResult[106] ? _T_2 : io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 194:16]
  wire [161:0] sigSum = {_T_3,io_mulAddResult[105:0],io_fromPreMul_bit0AlignedSigC}; // @[Cat.scala 29:58]
  wire [1:0] _T_6 = {1'b0,$signed(io_fromPreMul_doSubMags)}; // @[MulAddRecFN.scala 205:69]
  wire [12:0] _GEN_0 = {{11{_T_6[1]}},_T_6}; // @[MulAddRecFN.scala 205:43]
  wire [12:0] CDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_0); // @[MulAddRecFN.scala 205:43]
  wire [107:0] _T_10 = ~sigSum[161:54]; // @[MulAddRecFN.scala 208:13]
  wire [107:0] _T_14 = {1'h0,io_fromPreMul_highAlignedSigC[54:53],sigSum[159:55]}; // @[Cat.scala 29:58]
  wire [107:0] CDom_absSigSum = io_fromPreMul_doSubMags ? _T_10 : _T_14; // @[MulAddRecFN.scala 207:12]
  wire [52:0] _T_16 = ~sigSum[53:1]; // @[MulAddRecFN.scala 217:14]
  wire  _T_17 = |_T_16; // @[MulAddRecFN.scala 217:36]
  wire  _T_19 = |sigSum[54:1]; // @[MulAddRecFN.scala 218:37]
  wire  CDom_absSigSumExtra = io_fromPreMul_doSubMags ? _T_17 : _T_19; // @[MulAddRecFN.scala 216:12]
  wire [170:0] _GEN_1 = {{63'd0}, CDom_absSigSum}; // @[MulAddRecFN.scala 221:24]
  wire [170:0] _T_20 = _GEN_1 << io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 221:24]
  wire [57:0] CDom_mainSig = _T_20[107:50]; // @[MulAddRecFN.scala 221:56]
  wire [54:0] _T_22 = {CDom_absSigSum[52:0], 2'h0}; // @[MulAddRecFN.scala 224:53]
  wire  _T_25 = |_T_22[3:0]; // @[primitives.scala 121:54]
  wire  _T_27 = |_T_22[7:4]; // @[primitives.scala 121:54]
  wire  _T_29 = |_T_22[11:8]; // @[primitives.scala 121:54]
  wire  _T_31 = |_T_22[15:12]; // @[primitives.scala 121:54]
  wire  _T_33 = |_T_22[19:16]; // @[primitives.scala 121:54]
  wire  _T_35 = |_T_22[23:20]; // @[primitives.scala 121:54]
  wire  _T_37 = |_T_22[27:24]; // @[primitives.scala 121:54]
  wire  _T_39 = |_T_22[31:28]; // @[primitives.scala 121:54]
  wire  _T_41 = |_T_22[35:32]; // @[primitives.scala 121:54]
  wire  _T_43 = |_T_22[39:36]; // @[primitives.scala 121:54]
  wire  _T_45 = |_T_22[43:40]; // @[primitives.scala 121:54]
  wire  _T_47 = |_T_22[47:44]; // @[primitives.scala 121:54]
  wire  _T_49 = |_T_22[51:48]; // @[primitives.scala 121:54]
  wire  _T_51 = |_T_22[54:52]; // @[primitives.scala 124:57]
  wire [6:0] _T_57 = {_T_37,_T_35,_T_33,_T_31,_T_29,_T_27,_T_25}; // @[primitives.scala 125:20]
  wire [13:0] _T_64 = {_T_51,_T_49,_T_47,_T_45,_T_43,_T_41,_T_39,_T_57}; // @[primitives.scala 125:20]
  wire [3:0] _T_66 = ~io_fromPreMul_CDom_CAlignDist[5:2]; // @[primitives.scala 51:21]
  wire [16:0] _T_67 = -17'sh10000 >>> _T_66; // @[primitives.scala 77:58]
  wire [7:0] _T_73 = {{4'd0}, _T_67[8:5]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_75 = {_T_67[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_77 = _T_75 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_78 = _T_73 | _T_77; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_2 = {{2'd0}, _T_78[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_83 = _GEN_2 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_85 = {_T_78[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_87 = _T_85 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_88 = _T_83 | _T_87; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_3 = {{1'd0}, _T_88[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_93 = _GEN_3 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_95 = {_T_88[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_97 = _T_95 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_98 = _T_93 | _T_97; // @[Bitwise.scala 103:39]
  wire [12:0] _T_112 = {_T_98,_T_67[9],_T_67[10],_T_67[11],_T_67[12],_T_67[13]}; // @[Cat.scala 29:58]
  wire [13:0] _GEN_4 = {{1'd0}, _T_112}; // @[MulAddRecFN.scala 224:72]
  wire [13:0] _T_113 = _T_64 & _GEN_4; // @[MulAddRecFN.scala 224:72]
  wire  CDom_reduced4SigExtra = |_T_113; // @[MulAddRecFN.scala 225:73]
  wire  _T_116 = |CDom_mainSig[2:0]; // @[MulAddRecFN.scala 228:32]
  wire  _T_117 = _T_116 | CDom_reduced4SigExtra; // @[MulAddRecFN.scala 228:36]
  wire  _T_118 = _T_117 | CDom_absSigSumExtra; // @[MulAddRecFN.scala 228:61]
  wire [55:0] CDom_sig = {CDom_mainSig[57:3],_T_118}; // @[Cat.scala 29:58]
  wire  notCDom_signSigSum = sigSum[109]; // @[MulAddRecFN.scala 234:36]
  wire [108:0] _T_120 = ~sigSum[108:0]; // @[MulAddRecFN.scala 237:13]
  wire [108:0] _GEN_5 = {{108'd0}, io_fromPreMul_doSubMags}; // @[MulAddRecFN.scala 238:41]
  wire [108:0] _T_123 = sigSum[108:0] + _GEN_5; // @[MulAddRecFN.scala 238:41]
  wire [108:0] notCDom_absSigSum = notCDom_signSigSum ? _T_120 : _T_123; // @[MulAddRecFN.scala 236:12]
  wire  _T_126 = |notCDom_absSigSum[1:0]; // @[primitives.scala 104:54]
  wire  _T_128 = |notCDom_absSigSum[3:2]; // @[primitives.scala 104:54]
  wire  _T_130 = |notCDom_absSigSum[5:4]; // @[primitives.scala 104:54]
  wire  _T_132 = |notCDom_absSigSum[7:6]; // @[primitives.scala 104:54]
  wire  _T_134 = |notCDom_absSigSum[9:8]; // @[primitives.scala 104:54]
  wire  _T_136 = |notCDom_absSigSum[11:10]; // @[primitives.scala 104:54]
  wire  _T_138 = |notCDom_absSigSum[13:12]; // @[primitives.scala 104:54]
  wire  _T_140 = |notCDom_absSigSum[15:14]; // @[primitives.scala 104:54]
  wire  _T_142 = |notCDom_absSigSum[17:16]; // @[primitives.scala 104:54]
  wire  _T_144 = |notCDom_absSigSum[19:18]; // @[primitives.scala 104:54]
  wire  _T_146 = |notCDom_absSigSum[21:20]; // @[primitives.scala 104:54]
  wire  _T_148 = |notCDom_absSigSum[23:22]; // @[primitives.scala 104:54]
  wire  _T_150 = |notCDom_absSigSum[25:24]; // @[primitives.scala 104:54]
  wire  _T_152 = |notCDom_absSigSum[27:26]; // @[primitives.scala 104:54]
  wire  _T_154 = |notCDom_absSigSum[29:28]; // @[primitives.scala 104:54]
  wire  _T_156 = |notCDom_absSigSum[31:30]; // @[primitives.scala 104:54]
  wire  _T_158 = |notCDom_absSigSum[33:32]; // @[primitives.scala 104:54]
  wire  _T_160 = |notCDom_absSigSum[35:34]; // @[primitives.scala 104:54]
  wire  _T_162 = |notCDom_absSigSum[37:36]; // @[primitives.scala 104:54]
  wire  _T_164 = |notCDom_absSigSum[39:38]; // @[primitives.scala 104:54]
  wire  _T_166 = |notCDom_absSigSum[41:40]; // @[primitives.scala 104:54]
  wire  _T_168 = |notCDom_absSigSum[43:42]; // @[primitives.scala 104:54]
  wire  _T_170 = |notCDom_absSigSum[45:44]; // @[primitives.scala 104:54]
  wire  _T_172 = |notCDom_absSigSum[47:46]; // @[primitives.scala 104:54]
  wire  _T_174 = |notCDom_absSigSum[49:48]; // @[primitives.scala 104:54]
  wire  _T_176 = |notCDom_absSigSum[51:50]; // @[primitives.scala 104:54]
  wire  _T_178 = |notCDom_absSigSum[53:52]; // @[primitives.scala 104:54]
  wire  _T_180 = |notCDom_absSigSum[55:54]; // @[primitives.scala 104:54]
  wire  _T_182 = |notCDom_absSigSum[57:56]; // @[primitives.scala 104:54]
  wire  _T_184 = |notCDom_absSigSum[59:58]; // @[primitives.scala 104:54]
  wire  _T_186 = |notCDom_absSigSum[61:60]; // @[primitives.scala 104:54]
  wire  _T_188 = |notCDom_absSigSum[63:62]; // @[primitives.scala 104:54]
  wire  _T_190 = |notCDom_absSigSum[65:64]; // @[primitives.scala 104:54]
  wire  _T_192 = |notCDom_absSigSum[67:66]; // @[primitives.scala 104:54]
  wire  _T_194 = |notCDom_absSigSum[69:68]; // @[primitives.scala 104:54]
  wire  _T_196 = |notCDom_absSigSum[71:70]; // @[primitives.scala 104:54]
  wire  _T_198 = |notCDom_absSigSum[73:72]; // @[primitives.scala 104:54]
  wire  _T_200 = |notCDom_absSigSum[75:74]; // @[primitives.scala 104:54]
  wire  _T_202 = |notCDom_absSigSum[77:76]; // @[primitives.scala 104:54]
  wire  _T_204 = |notCDom_absSigSum[79:78]; // @[primitives.scala 104:54]
  wire  _T_206 = |notCDom_absSigSum[81:80]; // @[primitives.scala 104:54]
  wire  _T_208 = |notCDom_absSigSum[83:82]; // @[primitives.scala 104:54]
  wire  _T_210 = |notCDom_absSigSum[85:84]; // @[primitives.scala 104:54]
  wire  _T_212 = |notCDom_absSigSum[87:86]; // @[primitives.scala 104:54]
  wire  _T_214 = |notCDom_absSigSum[89:88]; // @[primitives.scala 104:54]
  wire  _T_216 = |notCDom_absSigSum[91:90]; // @[primitives.scala 104:54]
  wire  _T_218 = |notCDom_absSigSum[93:92]; // @[primitives.scala 104:54]
  wire  _T_220 = |notCDom_absSigSum[95:94]; // @[primitives.scala 104:54]
  wire  _T_222 = |notCDom_absSigSum[97:96]; // @[primitives.scala 104:54]
  wire  _T_224 = |notCDom_absSigSum[99:98]; // @[primitives.scala 104:54]
  wire  _T_226 = |notCDom_absSigSum[101:100]; // @[primitives.scala 104:54]
  wire  _T_228 = |notCDom_absSigSum[103:102]; // @[primitives.scala 104:54]
  wire  _T_230 = |notCDom_absSigSum[105:104]; // @[primitives.scala 104:54]
  wire  _T_232 = |notCDom_absSigSum[107:106]; // @[primitives.scala 104:54]
  wire  _T_234 = |notCDom_absSigSum[108]; // @[primitives.scala 107:57]
  wire [5:0] _T_239 = {_T_136,_T_134,_T_132,_T_130,_T_128,_T_126}; // @[primitives.scala 108:20]
  wire [12:0] _T_246 = {_T_150,_T_148,_T_146,_T_144,_T_142,_T_140,_T_138,_T_239}; // @[primitives.scala 108:20]
  wire [6:0] _T_252 = {_T_164,_T_162,_T_160,_T_158,_T_156,_T_154,_T_152}; // @[primitives.scala 108:20]
  wire [26:0] _T_260 = {_T_178,_T_176,_T_174,_T_172,_T_170,_T_168,_T_166,_T_252,_T_246}; // @[primitives.scala 108:20]
  wire [6:0] _T_266 = {_T_192,_T_190,_T_188,_T_186,_T_184,_T_182,_T_180}; // @[primitives.scala 108:20]
  wire [13:0] _T_273 = {_T_206,_T_204,_T_202,_T_200,_T_198,_T_196,_T_194,_T_266}; // @[primitives.scala 108:20]
  wire [6:0] _T_279 = {_T_220,_T_218,_T_216,_T_214,_T_212,_T_210,_T_208}; // @[primitives.scala 108:20]
  wire [54:0] notCDom_reduced2AbsSigSum = {_T_234,_T_232,_T_230,_T_228,_T_226,_T_224,_T_222,_T_279,_T_273,_T_260}; // @[primitives.scala 108:20]
  wire [5:0] _T_343 = notCDom_reduced2AbsSigSum[1] ? 6'h35 : 6'h36; // @[Mux.scala 47:69]
  wire [5:0] _T_344 = notCDom_reduced2AbsSigSum[2] ? 6'h34 : _T_343; // @[Mux.scala 47:69]
  wire [5:0] _T_345 = notCDom_reduced2AbsSigSum[3] ? 6'h33 : _T_344; // @[Mux.scala 47:69]
  wire [5:0] _T_346 = notCDom_reduced2AbsSigSum[4] ? 6'h32 : _T_345; // @[Mux.scala 47:69]
  wire [5:0] _T_347 = notCDom_reduced2AbsSigSum[5] ? 6'h31 : _T_346; // @[Mux.scala 47:69]
  wire [5:0] _T_348 = notCDom_reduced2AbsSigSum[6] ? 6'h30 : _T_347; // @[Mux.scala 47:69]
  wire [5:0] _T_349 = notCDom_reduced2AbsSigSum[7] ? 6'h2f : _T_348; // @[Mux.scala 47:69]
  wire [5:0] _T_350 = notCDom_reduced2AbsSigSum[8] ? 6'h2e : _T_349; // @[Mux.scala 47:69]
  wire [5:0] _T_351 = notCDom_reduced2AbsSigSum[9] ? 6'h2d : _T_350; // @[Mux.scala 47:69]
  wire [5:0] _T_352 = notCDom_reduced2AbsSigSum[10] ? 6'h2c : _T_351; // @[Mux.scala 47:69]
  wire [5:0] _T_353 = notCDom_reduced2AbsSigSum[11] ? 6'h2b : _T_352; // @[Mux.scala 47:69]
  wire [5:0] _T_354 = notCDom_reduced2AbsSigSum[12] ? 6'h2a : _T_353; // @[Mux.scala 47:69]
  wire [5:0] _T_355 = notCDom_reduced2AbsSigSum[13] ? 6'h29 : _T_354; // @[Mux.scala 47:69]
  wire [5:0] _T_356 = notCDom_reduced2AbsSigSum[14] ? 6'h28 : _T_355; // @[Mux.scala 47:69]
  wire [5:0] _T_357 = notCDom_reduced2AbsSigSum[15] ? 6'h27 : _T_356; // @[Mux.scala 47:69]
  wire [5:0] _T_358 = notCDom_reduced2AbsSigSum[16] ? 6'h26 : _T_357; // @[Mux.scala 47:69]
  wire [5:0] _T_359 = notCDom_reduced2AbsSigSum[17] ? 6'h25 : _T_358; // @[Mux.scala 47:69]
  wire [5:0] _T_360 = notCDom_reduced2AbsSigSum[18] ? 6'h24 : _T_359; // @[Mux.scala 47:69]
  wire [5:0] _T_361 = notCDom_reduced2AbsSigSum[19] ? 6'h23 : _T_360; // @[Mux.scala 47:69]
  wire [5:0] _T_362 = notCDom_reduced2AbsSigSum[20] ? 6'h22 : _T_361; // @[Mux.scala 47:69]
  wire [5:0] _T_363 = notCDom_reduced2AbsSigSum[21] ? 6'h21 : _T_362; // @[Mux.scala 47:69]
  wire [5:0] _T_364 = notCDom_reduced2AbsSigSum[22] ? 6'h20 : _T_363; // @[Mux.scala 47:69]
  wire [5:0] _T_365 = notCDom_reduced2AbsSigSum[23] ? 6'h1f : _T_364; // @[Mux.scala 47:69]
  wire [5:0] _T_366 = notCDom_reduced2AbsSigSum[24] ? 6'h1e : _T_365; // @[Mux.scala 47:69]
  wire [5:0] _T_367 = notCDom_reduced2AbsSigSum[25] ? 6'h1d : _T_366; // @[Mux.scala 47:69]
  wire [5:0] _T_368 = notCDom_reduced2AbsSigSum[26] ? 6'h1c : _T_367; // @[Mux.scala 47:69]
  wire [5:0] _T_369 = notCDom_reduced2AbsSigSum[27] ? 6'h1b : _T_368; // @[Mux.scala 47:69]
  wire [5:0] _T_370 = notCDom_reduced2AbsSigSum[28] ? 6'h1a : _T_369; // @[Mux.scala 47:69]
  wire [5:0] _T_371 = notCDom_reduced2AbsSigSum[29] ? 6'h19 : _T_370; // @[Mux.scala 47:69]
  wire [5:0] _T_372 = notCDom_reduced2AbsSigSum[30] ? 6'h18 : _T_371; // @[Mux.scala 47:69]
  wire [5:0] _T_373 = notCDom_reduced2AbsSigSum[31] ? 6'h17 : _T_372; // @[Mux.scala 47:69]
  wire [5:0] _T_374 = notCDom_reduced2AbsSigSum[32] ? 6'h16 : _T_373; // @[Mux.scala 47:69]
  wire [5:0] _T_375 = notCDom_reduced2AbsSigSum[33] ? 6'h15 : _T_374; // @[Mux.scala 47:69]
  wire [5:0] _T_376 = notCDom_reduced2AbsSigSum[34] ? 6'h14 : _T_375; // @[Mux.scala 47:69]
  wire [5:0] _T_377 = notCDom_reduced2AbsSigSum[35] ? 6'h13 : _T_376; // @[Mux.scala 47:69]
  wire [5:0] _T_378 = notCDom_reduced2AbsSigSum[36] ? 6'h12 : _T_377; // @[Mux.scala 47:69]
  wire [5:0] _T_379 = notCDom_reduced2AbsSigSum[37] ? 6'h11 : _T_378; // @[Mux.scala 47:69]
  wire [5:0] _T_380 = notCDom_reduced2AbsSigSum[38] ? 6'h10 : _T_379; // @[Mux.scala 47:69]
  wire [5:0] _T_381 = notCDom_reduced2AbsSigSum[39] ? 6'hf : _T_380; // @[Mux.scala 47:69]
  wire [5:0] _T_382 = notCDom_reduced2AbsSigSum[40] ? 6'he : _T_381; // @[Mux.scala 47:69]
  wire [5:0] _T_383 = notCDom_reduced2AbsSigSum[41] ? 6'hd : _T_382; // @[Mux.scala 47:69]
  wire [5:0] _T_384 = notCDom_reduced2AbsSigSum[42] ? 6'hc : _T_383; // @[Mux.scala 47:69]
  wire [5:0] _T_385 = notCDom_reduced2AbsSigSum[43] ? 6'hb : _T_384; // @[Mux.scala 47:69]
  wire [5:0] _T_386 = notCDom_reduced2AbsSigSum[44] ? 6'ha : _T_385; // @[Mux.scala 47:69]
  wire [5:0] _T_387 = notCDom_reduced2AbsSigSum[45] ? 6'h9 : _T_386; // @[Mux.scala 47:69]
  wire [5:0] _T_388 = notCDom_reduced2AbsSigSum[46] ? 6'h8 : _T_387; // @[Mux.scala 47:69]
  wire [5:0] _T_389 = notCDom_reduced2AbsSigSum[47] ? 6'h7 : _T_388; // @[Mux.scala 47:69]
  wire [5:0] _T_390 = notCDom_reduced2AbsSigSum[48] ? 6'h6 : _T_389; // @[Mux.scala 47:69]
  wire [5:0] _T_391 = notCDom_reduced2AbsSigSum[49] ? 6'h5 : _T_390; // @[Mux.scala 47:69]
  wire [5:0] _T_392 = notCDom_reduced2AbsSigSum[50] ? 6'h4 : _T_391; // @[Mux.scala 47:69]
  wire [5:0] _T_393 = notCDom_reduced2AbsSigSum[51] ? 6'h3 : _T_392; // @[Mux.scala 47:69]
  wire [5:0] _T_394 = notCDom_reduced2AbsSigSum[52] ? 6'h2 : _T_393; // @[Mux.scala 47:69]
  wire [5:0] _T_395 = notCDom_reduced2AbsSigSum[53] ? 6'h1 : _T_394; // @[Mux.scala 47:69]
  wire [5:0] notCDom_normDistReduced2 = notCDom_reduced2AbsSigSum[54] ? 6'h0 : _T_395; // @[Mux.scala 47:69]
  wire [6:0] notCDom_nearNormDist = {notCDom_normDistReduced2, 1'h0}; // @[MulAddRecFN.scala 242:56]
  wire [7:0] _T_396 = {1'b0,$signed(notCDom_nearNormDist)}; // @[MulAddRecFN.scala 243:69]
  wire [12:0] _GEN_6 = {{5{_T_396[7]}},_T_396}; // @[MulAddRecFN.scala 243:46]
  wire [12:0] notCDom_sExp = $signed(io_fromPreMul_sExpSum) - $signed(_GEN_6); // @[MulAddRecFN.scala 243:46]
  wire [235:0] _GEN_7 = {{127'd0}, notCDom_absSigSum}; // @[MulAddRecFN.scala 245:27]
  wire [235:0] _T_399 = _GEN_7 << notCDom_nearNormDist; // @[MulAddRecFN.scala 245:27]
  wire [57:0] notCDom_mainSig = _T_399[109:52]; // @[MulAddRecFN.scala 245:50]
  wire  _T_404 = |notCDom_reduced2AbsSigSum[1:0]; // @[primitives.scala 104:54]
  wire  _T_406 = |notCDom_reduced2AbsSigSum[3:2]; // @[primitives.scala 104:54]
  wire  _T_408 = |notCDom_reduced2AbsSigSum[5:4]; // @[primitives.scala 104:54]
  wire  _T_410 = |notCDom_reduced2AbsSigSum[7:6]; // @[primitives.scala 104:54]
  wire  _T_412 = |notCDom_reduced2AbsSigSum[9:8]; // @[primitives.scala 104:54]
  wire  _T_414 = |notCDom_reduced2AbsSigSum[11:10]; // @[primitives.scala 104:54]
  wire  _T_416 = |notCDom_reduced2AbsSigSum[13:12]; // @[primitives.scala 104:54]
  wire  _T_418 = |notCDom_reduced2AbsSigSum[15:14]; // @[primitives.scala 104:54]
  wire  _T_420 = |notCDom_reduced2AbsSigSum[17:16]; // @[primitives.scala 104:54]
  wire  _T_422 = |notCDom_reduced2AbsSigSum[19:18]; // @[primitives.scala 104:54]
  wire  _T_424 = |notCDom_reduced2AbsSigSum[21:20]; // @[primitives.scala 104:54]
  wire  _T_426 = |notCDom_reduced2AbsSigSum[23:22]; // @[primitives.scala 104:54]
  wire  _T_428 = |notCDom_reduced2AbsSigSum[25:24]; // @[primitives.scala 104:54]
  wire  _T_430 = |notCDom_reduced2AbsSigSum[26]; // @[primitives.scala 107:57]
  wire [6:0] _T_436 = {_T_416,_T_414,_T_412,_T_410,_T_408,_T_406,_T_404}; // @[primitives.scala 108:20]
  wire [13:0] _T_443 = {_T_430,_T_428,_T_426,_T_424,_T_422,_T_420,_T_418,_T_436}; // @[primitives.scala 108:20]
  wire [4:0] _T_445 = ~notCDom_normDistReduced2[5:1]; // @[primitives.scala 51:21]
  wire [32:0] _T_446 = -33'sh100000000 >>> _T_445; // @[primitives.scala 77:58]
  wire [7:0] _T_452 = {{4'd0}, _T_446[8:5]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_454 = {_T_446[4:1], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_456 = _T_454 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_457 = _T_452 | _T_456; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_8 = {{2'd0}, _T_457[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_462 = _GEN_8 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_464 = {_T_457[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_466 = _T_464 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_467 = _T_462 | _T_466; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_9 = {{1'd0}, _T_467[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_472 = _GEN_9 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_474 = {_T_467[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_476 = _T_474 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_477 = _T_472 | _T_476; // @[Bitwise.scala 103:39]
  wire [12:0] _T_491 = {_T_477,_T_446[9],_T_446[10],_T_446[11],_T_446[12],_T_446[13]}; // @[Cat.scala 29:58]
  wire [13:0] _GEN_10 = {{1'd0}, _T_491}; // @[MulAddRecFN.scala 249:78]
  wire [13:0] _T_492 = _T_443 & _GEN_10; // @[MulAddRecFN.scala 249:78]
  wire  notCDom_reduced4SigExtra = |_T_492; // @[MulAddRecFN.scala 251:11]
  wire  _T_495 = |notCDom_mainSig[2:0]; // @[MulAddRecFN.scala 254:35]
  wire  _T_496 = _T_495 | notCDom_reduced4SigExtra; // @[MulAddRecFN.scala 254:39]
  wire [55:0] notCDom_sig = {notCDom_mainSig[57:3],_T_496}; // @[Cat.scala 29:58]
  wire  notCDom_completeCancellation = notCDom_sig[55:54] == 2'h0; // @[MulAddRecFN.scala 257:50]
  wire  _T_498 = io_fromPreMul_signProd ^ notCDom_signSigSum; // @[MulAddRecFN.scala 261:36]
  wire  notCDom_sign = notCDom_completeCancellation ? 1'h0 : _T_498; // @[MulAddRecFN.scala 259:12]
  wire  notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB; // @[MulAddRecFN.scala 266:49]
  wire  notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 267:44]
  wire  _T_499 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 269:32]
  wire  notNaN_addZeros = _T_499 & io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 269:58]
  wire  _T_500 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 274:31]
  wire  _T_501 = io_fromPreMul_isSigNaNAny | _T_500; // @[MulAddRecFN.scala 273:35]
  wire  _T_502 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB; // @[MulAddRecFN.scala 275:32]
  wire  _T_503 = _T_501 | _T_502; // @[MulAddRecFN.scala 274:57]
  wire  _T_504 = ~io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 276:10]
  wire  _T_506 = _T_504 & notNaN_isInfProd; // @[MulAddRecFN.scala 276:36]
  wire  _T_507 = _T_506 & io_fromPreMul_isInfC; // @[MulAddRecFN.scala 277:61]
  wire  _T_508 = _T_507 & io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 278:35]
  wire  _T_511 = ~io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 285:14]
  wire  _T_512 = _T_511 & notCDom_completeCancellation; // @[MulAddRecFN.scala 285:42]
  wire  _T_514 = notNaN_isInfProd & io_fromPreMul_signProd; // @[MulAddRecFN.scala 287:27]
  wire  _T_515 = io_fromPreMul_isInfC & CDom_sign; // @[MulAddRecFN.scala 288:31]
  wire  _T_516 = _T_514 | _T_515; // @[MulAddRecFN.scala 287:54]
  wire  _T_519 = notNaN_addZeros & io_fromPreMul_signProd; // @[MulAddRecFN.scala 289:48]
  wire  _T_520 = _T_519 & CDom_sign; // @[MulAddRecFN.scala 290:36]
  wire  _T_521 = _T_516 | _T_520; // @[MulAddRecFN.scala 288:43]
  wire  _T_526 = ~notNaN_isInfOut; // @[MulAddRecFN.scala 293:10]
  wire  _T_527 = ~notNaN_addZeros; // @[MulAddRecFN.scala 293:31]
  wire  _T_528 = _T_526 & _T_527; // @[MulAddRecFN.scala 293:28]
  wire  _T_529 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign; // @[MulAddRecFN.scala 294:17]
  wire  _T_530 = _T_528 & _T_529; // @[MulAddRecFN.scala 293:49]
  assign io_invalidExc = _T_503 | _T_508; // @[MulAddRecFN.scala 272:19]
  assign io_rawOut_isNaN = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 280:21]
  assign io_rawOut_isInf = notNaN_isInfProd | io_fromPreMul_isInfC; // @[MulAddRecFN.scala 281:21]
  assign io_rawOut_isZero = notNaN_addZeros | _T_512; // @[MulAddRecFN.scala 283:22]
  assign io_rawOut_sign = _T_521 | _T_530; // @[MulAddRecFN.scala 286:20]
  assign io_rawOut_sExp = io_fromPreMul_CIsDominant ? $signed(CDom_sExp) : $signed(notCDom_sExp); // @[MulAddRecFN.scala 295:20]
  assign io_rawOut_sig = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig; // @[MulAddRecFN.scala 296:19]
endmodule
module RoundAnyRawFNToRecFN_2(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  output [64:0] io_out
);
  wire  doShiftSigDown1 = io_in_sig[55]; // @[RoundAnyRawFNToRecFN.scala 118:61]
  wire [11:0] _T_4 = ~io_in_sExp[11:0]; // @[primitives.scala 51:21]
  wire [64:0] _T_17 = -65'sh10000000000000000 >>> _T_4[5:0]; // @[primitives.scala 77:58]
  wire [31:0] _T_23 = {{16'd0}, _T_17[44:29]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_25 = {_T_17[28:13], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_27 = _T_25 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_28 = _T_23 | _T_27; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _T_28[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_33 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_35 = {_T_28[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_37 = _T_35 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_38 = _T_33 | _T_37; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _T_38[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_43 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_45 = {_T_38[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_47 = _T_45 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_48 = _T_43 | _T_47; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _T_48[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_53 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_55 = {_T_48[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_57 = _T_55 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_58 = _T_53 | _T_57; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _T_58[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_63 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_65 = {_T_58[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_67 = _T_65 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_68 = _T_63 | _T_67; // @[Bitwise.scala 103:39]
  wire [15:0] _T_74 = {{8'd0}, _T_17[60:53]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_76 = {_T_17[52:45], 8'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_78 = _T_76 & 16'hff00; // @[Bitwise.scala 103:75]
  wire [15:0] _T_79 = _T_74 | _T_78; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_4 = {{4'd0}, _T_79[15:4]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_84 = _GEN_4 & 16'hf0f; // @[Bitwise.scala 103:31]
  wire [15:0] _T_86 = {_T_79[11:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_88 = _T_86 & 16'hf0f0; // @[Bitwise.scala 103:75]
  wire [15:0] _T_89 = _T_84 | _T_88; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_5 = {{2'd0}, _T_89[15:2]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_94 = _GEN_5 & 16'h3333; // @[Bitwise.scala 103:31]
  wire [15:0] _T_96 = {_T_89[13:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_98 = _T_96 & 16'hcccc; // @[Bitwise.scala 103:75]
  wire [15:0] _T_99 = _T_94 | _T_98; // @[Bitwise.scala 103:39]
  wire [15:0] _GEN_6 = {{1'd0}, _T_99[15:1]}; // @[Bitwise.scala 103:31]
  wire [15:0] _T_104 = _GEN_6 & 16'h5555; // @[Bitwise.scala 103:31]
  wire [15:0] _T_106 = {_T_99[14:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [15:0] _T_108 = _T_106 & 16'haaaa; // @[Bitwise.scala 103:75]
  wire [15:0] _T_109 = _T_104 | _T_108; // @[Bitwise.scala 103:39]
  wire [50:0] _T_118 = {_T_68,_T_109,_T_17[61],_T_17[62],_T_17[63]}; // @[Cat.scala 29:58]
  wire [50:0] _T_119 = ~_T_118; // @[primitives.scala 74:36]
  wire [50:0] _T_120 = _T_4[6] ? 51'h0 : _T_119; // @[primitives.scala 74:21]
  wire [50:0] _T_121 = ~_T_120; // @[primitives.scala 74:17]
  wire [50:0] _T_122 = ~_T_121; // @[primitives.scala 74:36]
  wire [50:0] _T_123 = _T_4[7] ? 51'h0 : _T_122; // @[primitives.scala 74:21]
  wire [50:0] _T_124 = ~_T_123; // @[primitives.scala 74:17]
  wire [50:0] _T_125 = ~_T_124; // @[primitives.scala 74:36]
  wire [50:0] _T_126 = _T_4[8] ? 51'h0 : _T_125; // @[primitives.scala 74:21]
  wire [50:0] _T_127 = ~_T_126; // @[primitives.scala 74:17]
  wire [50:0] _T_128 = ~_T_127; // @[primitives.scala 74:36]
  wire [50:0] _T_129 = _T_4[9] ? 51'h0 : _T_128; // @[primitives.scala 74:21]
  wire [50:0] _T_130 = ~_T_129; // @[primitives.scala 74:17]
  wire [53:0] _T_131 = {_T_130,3'h7}; // @[Cat.scala 29:58]
  wire [2:0] _T_147 = {_T_17[0],_T_17[1],_T_17[2]}; // @[Cat.scala 29:58]
  wire [2:0] _T_148 = _T_4[6] ? _T_147 : 3'h0; // @[primitives.scala 61:24]
  wire [2:0] _T_149 = _T_4[7] ? _T_148 : 3'h0; // @[primitives.scala 61:24]
  wire [2:0] _T_150 = _T_4[8] ? _T_149 : 3'h0; // @[primitives.scala 61:24]
  wire [2:0] _T_151 = _T_4[9] ? _T_150 : 3'h0; // @[primitives.scala 61:24]
  wire [53:0] _T_152 = _T_4[10] ? _T_131 : {{51'd0}, _T_151}; // @[primitives.scala 66:24]
  wire [53:0] _T_153 = _T_4[11] ? _T_152 : 54'h0; // @[primitives.scala 61:24]
  wire [53:0] _GEN_7 = {{53'd0}, doShiftSigDown1}; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [53:0] _T_154 = _T_153 | _GEN_7; // @[RoundAnyRawFNToRecFN.scala 157:23]
  wire [55:0] _T_155 = {_T_154,2'h3}; // @[Cat.scala 29:58]
  wire [55:0] _T_157 = {1'h0,_T_155[55:1]}; // @[Cat.scala 29:58]
  wire [55:0] _T_158 = ~_T_157; // @[RoundAnyRawFNToRecFN.scala 161:28]
  wire [55:0] _T_159 = _T_158 & _T_155; // @[RoundAnyRawFNToRecFN.scala 161:46]
  wire [55:0] _T_160 = io_in_sig & _T_159; // @[RoundAnyRawFNToRecFN.scala 162:40]
  wire  _T_161 = |_T_160; // @[RoundAnyRawFNToRecFN.scala 162:56]
  wire [55:0] _T_162 = io_in_sig & _T_157; // @[RoundAnyRawFNToRecFN.scala 163:42]
  wire  _T_163 = |_T_162; // @[RoundAnyRawFNToRecFN.scala 163:62]
  wire  _T_164 = _T_161 | _T_163; // @[RoundAnyRawFNToRecFN.scala 164:36]
  wire [55:0] _T_179 = ~_T_155; // @[RoundAnyRawFNToRecFN.scala 178:32]
  wire [55:0] _T_180 = io_in_sig & _T_179; // @[RoundAnyRawFNToRecFN.scala 178:30]
  wire [54:0] _T_184 = _T_164 ? _T_159[55:1] : 55'h0; // @[RoundAnyRawFNToRecFN.scala 179:24]
  wire [54:0] _GEN_8 = {{1'd0}, _T_180[55:2]}; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [54:0] _T_185 = _GEN_8 | _T_184; // @[RoundAnyRawFNToRecFN.scala 178:47]
  wire [2:0] _T_188 = {1'b0,$signed(_T_185[54:53])}; // @[RoundAnyRawFNToRecFN.scala 183:69]
  wire [12:0] _GEN_9 = {{10{_T_188[2]}},_T_188}; // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [13:0] _T_189 = $signed(io_in_sExp) + $signed(_GEN_9); // @[RoundAnyRawFNToRecFN.scala 183:40]
  wire [11:0] common_expOut = _T_189[11:0]; // @[RoundAnyRawFNToRecFN.scala 185:37]
  wire [51:0] common_fractOut = doShiftSigDown1 ? _T_185[52:1] : _T_185[51:0]; // @[RoundAnyRawFNToRecFN.scala 187:16]
  wire [3:0] _T_194 = _T_189[13:10]; // @[RoundAnyRawFNToRecFN.scala 194:30]
  wire  common_overflow = $signed(_T_194) >= 4'sh3; // @[RoundAnyRawFNToRecFN.scala 194:50]
  wire  common_totalUnderflow = $signed(_T_189) < 14'sh3ce; // @[RoundAnyRawFNToRecFN.scala 198:31]
  wire  isNaNOut = io_invalidExc | io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 233:34]
  wire  _T_232 = ~isNaNOut; // @[RoundAnyRawFNToRecFN.scala 235:22]
  wire  _T_233 = ~io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 235:36]
  wire  _T_234 = _T_232 & _T_233; // @[RoundAnyRawFNToRecFN.scala 235:33]
  wire  _T_235 = ~io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 235:64]
  wire  commonCase = _T_234 & _T_235; // @[RoundAnyRawFNToRecFN.scala 235:61]
  wire  overflow = commonCase & common_overflow; // @[RoundAnyRawFNToRecFN.scala 236:32]
  wire  pegMinNonzeroMagOut = commonCase & common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 243:20]
  wire  signOut = isNaNOut ? 1'h0 : io_in_sign; // @[RoundAnyRawFNToRecFN.scala 248:22]
  wire  _T_242 = io_in_isZero | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 251:32]
  wire [11:0] _T_243 = _T_242 ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 251:18]
  wire [11:0] _T_244 = ~_T_243; // @[RoundAnyRawFNToRecFN.scala 251:14]
  wire [11:0] _T_245 = common_expOut & _T_244; // @[RoundAnyRawFNToRecFN.scala 250:24]
  wire [11:0] _T_247 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 255:18]
  wire [11:0] _T_248 = ~_T_247; // @[RoundAnyRawFNToRecFN.scala 255:14]
  wire [11:0] _T_249 = _T_245 & _T_248; // @[RoundAnyRawFNToRecFN.scala 254:17]
  wire [11:0] _T_250 = overflow ? 12'h400 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 259:18]
  wire [11:0] _T_251 = ~_T_250; // @[RoundAnyRawFNToRecFN.scala 259:14]
  wire [11:0] _T_252 = _T_249 & _T_251; // @[RoundAnyRawFNToRecFN.scala 258:17]
  wire [11:0] _T_253 = io_in_isInf ? 12'h200 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 263:18]
  wire [11:0] _T_254 = ~_T_253; // @[RoundAnyRawFNToRecFN.scala 263:14]
  wire [11:0] _T_255 = _T_252 & _T_254; // @[RoundAnyRawFNToRecFN.scala 262:17]
  wire [11:0] _T_256 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0; // @[RoundAnyRawFNToRecFN.scala 267:16]
  wire [11:0] _T_257 = _T_255 | _T_256; // @[RoundAnyRawFNToRecFN.scala 266:18]
  wire [11:0] _T_258 = overflow ? 12'hbff : 12'h0; // @[RoundAnyRawFNToRecFN.scala 271:16]
  wire [11:0] _T_259 = _T_257 | _T_258; // @[RoundAnyRawFNToRecFN.scala 270:15]
  wire [11:0] _T_260 = io_in_isInf ? 12'hc00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 275:16]
  wire [11:0] _T_261 = _T_259 | _T_260; // @[RoundAnyRawFNToRecFN.scala 274:15]
  wire [11:0] _T_262 = isNaNOut ? 12'he00 : 12'h0; // @[RoundAnyRawFNToRecFN.scala 276:16]
  wire [11:0] expOut = _T_261 | _T_262; // @[RoundAnyRawFNToRecFN.scala 275:77]
  wire  _T_263 = isNaNOut | io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 278:22]
  wire  _T_264 = _T_263 | common_totalUnderflow; // @[RoundAnyRawFNToRecFN.scala 278:38]
  wire [51:0] _T_265 = isNaNOut ? 52'h8000000000000 : 52'h0; // @[RoundAnyRawFNToRecFN.scala 279:16]
  wire [51:0] _T_266 = _T_264 ? _T_265 : common_fractOut; // @[RoundAnyRawFNToRecFN.scala 278:12]
  wire [51:0] _T_268 = overflow ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [51:0] fractOut = _T_266 | _T_268; // @[RoundAnyRawFNToRecFN.scala 281:11]
  wire [12:0] _T_269 = {signOut,expOut}; // @[Cat.scala 29:58]
  assign io_out = {_T_269,fractOut}; // @[RoundAnyRawFNToRecFN.scala 284:12]
endmodule
module RoundRawFNToRecFN(
  input         io_invalidExc,
  input         io_in_isNaN,
  input         io_in_isInf,
  input         io_in_isZero,
  input         io_in_sign,
  input  [12:0] io_in_sExp,
  input  [55:0] io_in_sig,
  output [64:0] io_out
);
  wire  roundAnyRawFNToRecFN_io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire  roundAnyRawFNToRecFN_io_in_sign; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [12:0] roundAnyRawFNToRecFN_io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [55:0] roundAnyRawFNToRecFN_io_in_sig; // @[RoundAnyRawFNToRecFN.scala 307:15]
  wire [64:0] roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 307:15]
  RoundAnyRawFNToRecFN_2 roundAnyRawFNToRecFN ( // @[RoundAnyRawFNToRecFN.scala 307:15]
    .io_invalidExc(roundAnyRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundAnyRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundAnyRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundAnyRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundAnyRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundAnyRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundAnyRawFNToRecFN_io_in_sig),
    .io_out(roundAnyRawFNToRecFN_io_out)
  );
  assign io_out = roundAnyRawFNToRecFN_io_out; // @[RoundAnyRawFNToRecFN.scala 315:23]
  assign roundAnyRawFNToRecFN_io_invalidExc = io_invalidExc; // @[RoundAnyRawFNToRecFN.scala 310:44]
  assign roundAnyRawFNToRecFN_io_in_isNaN = io_in_isNaN; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isInf = io_in_isInf; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_isZero = io_in_isZero; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sign = io_in_sign; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sExp = io_in_sExp; // @[RoundAnyRawFNToRecFN.scala 312:44]
  assign roundAnyRawFNToRecFN_io_in_sig = io_in_sig; // @[RoundAnyRawFNToRecFN.scala 312:44]
endmodule
module MulAddRecFN(
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  output [64:0] io_out
);
  wire [64:0] mulAddRecFNToRaw_preMul_io_a; // @[MulAddRecFN.scala 318:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_b; // @[MulAddRecFN.scala 318:15]
  wire [64:0] mulAddRecFNToRaw_preMul_io_c; // @[MulAddRecFN.scala 318:15]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddA; // @[MulAddRecFN.scala 318:15]
  wire [52:0] mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 318:15]
  wire [105:0] mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 318:15]
  wire [12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 318:15]
  wire [5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 318:15]
  wire [54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 318:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_signProd; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC; // @[MulAddRecFN.scala 320:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant; // @[MulAddRecFN.scala 320:15]
  wire [5:0] mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist; // @[MulAddRecFN.scala 320:15]
  wire [54:0] mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC; // @[MulAddRecFN.scala 320:15]
  wire [106:0] mulAddRecFNToRaw_postMul_io_mulAddResult; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 320:15]
  wire  mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 320:15]
  wire [12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 320:15]
  wire [55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 320:15]
  wire  roundRawFNToRecFN_io_invalidExc; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isNaN; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isInf; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_isZero; // @[MulAddRecFN.scala 340:15]
  wire  roundRawFNToRecFN_io_in_sign; // @[MulAddRecFN.scala 340:15]
  wire [12:0] roundRawFNToRecFN_io_in_sExp; // @[MulAddRecFN.scala 340:15]
  wire [55:0] roundRawFNToRecFN_io_in_sig; // @[MulAddRecFN.scala 340:15]
  wire [64:0] roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 340:15]
  wire [105:0] _T = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB; // @[MulAddRecFN.scala 328:45]
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul ( // @[MulAddRecFN.scala 318:15]
    .io_a(mulAddRecFNToRaw_preMul_io_a),
    .io_b(mulAddRecFNToRaw_preMul_io_b),
    .io_c(mulAddRecFNToRaw_preMul_io_c),
    .io_mulAddA(mulAddRecFNToRaw_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFNToRaw_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFNToRaw_preMul_io_mulAddC),
    .io_toPostMul_isSigNaNAny(mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny),
    .io_toPostMul_isNaNAOrB(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB),
    .io_toPostMul_isInfA(mulAddRecFNToRaw_preMul_io_toPostMul_isInfA),
    .io_toPostMul_isZeroA(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA),
    .io_toPostMul_isInfB(mulAddRecFNToRaw_preMul_io_toPostMul_isInfB),
    .io_toPostMul_isZeroB(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB),
    .io_toPostMul_signProd(mulAddRecFNToRaw_preMul_io_toPostMul_signProd),
    .io_toPostMul_isNaNC(mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC),
    .io_toPostMul_isInfC(mulAddRecFNToRaw_preMul_io_toPostMul_isInfC),
    .io_toPostMul_isZeroC(mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC),
    .io_toPostMul_sExpSum(mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_doSubMags(mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags),
    .io_toPostMul_CIsDominant(mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant),
    .io_toPostMul_CDom_CAlignDist(mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist),
    .io_toPostMul_highAlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC),
    .io_toPostMul_bit0AlignedSigC(mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC)
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul ( // @[MulAddRecFN.scala 320:15]
    .io_fromPreMul_isSigNaNAny(mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny),
    .io_fromPreMul_isNaNAOrB(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB),
    .io_fromPreMul_isInfA(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA),
    .io_fromPreMul_isZeroA(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA),
    .io_fromPreMul_isInfB(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB),
    .io_fromPreMul_isZeroB(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB),
    .io_fromPreMul_signProd(mulAddRecFNToRaw_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isNaNC(mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC),
    .io_fromPreMul_isInfC(mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC),
    .io_fromPreMul_isZeroC(mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC),
    .io_fromPreMul_sExpSum(mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_doSubMags(mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags),
    .io_fromPreMul_CIsDominant(mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant),
    .io_fromPreMul_CDom_CAlignDist(mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist),
    .io_fromPreMul_highAlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC),
    .io_fromPreMul_bit0AlignedSigC(mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC),
    .io_mulAddResult(mulAddRecFNToRaw_postMul_io_mulAddResult),
    .io_invalidExc(mulAddRecFNToRaw_postMul_io_invalidExc),
    .io_rawOut_isNaN(mulAddRecFNToRaw_postMul_io_rawOut_isNaN),
    .io_rawOut_isInf(mulAddRecFNToRaw_postMul_io_rawOut_isInf),
    .io_rawOut_isZero(mulAddRecFNToRaw_postMul_io_rawOut_isZero),
    .io_rawOut_sign(mulAddRecFNToRaw_postMul_io_rawOut_sign),
    .io_rawOut_sExp(mulAddRecFNToRaw_postMul_io_rawOut_sExp),
    .io_rawOut_sig(mulAddRecFNToRaw_postMul_io_rawOut_sig)
  );
  RoundRawFNToRecFN roundRawFNToRecFN ( // @[MulAddRecFN.scala 340:15]
    .io_invalidExc(roundRawFNToRecFN_io_invalidExc),
    .io_in_isNaN(roundRawFNToRecFN_io_in_isNaN),
    .io_in_isInf(roundRawFNToRecFN_io_in_isInf),
    .io_in_isZero(roundRawFNToRecFN_io_in_isZero),
    .io_in_sign(roundRawFNToRecFN_io_in_sign),
    .io_in_sExp(roundRawFNToRecFN_io_in_sExp),
    .io_in_sig(roundRawFNToRecFN_io_in_sig),
    .io_out(roundRawFNToRecFN_io_out)
  );
  assign io_out = roundRawFNToRecFN_io_out; // @[MulAddRecFN.scala 346:23]
  assign mulAddRecFNToRaw_preMul_io_a = io_a; // @[MulAddRecFN.scala 323:35]
  assign mulAddRecFNToRaw_preMul_io_b = io_b; // @[MulAddRecFN.scala 324:35]
  assign mulAddRecFNToRaw_preMul_io_c = io_c; // @[MulAddRecFN.scala 325:35]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isSigNaNAny = mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNAOrB = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfA = mulAddRecFNToRaw_preMul_io_toPostMul_isInfA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroA = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfB = mulAddRecFNToRaw_preMul_io_toPostMul_isInfB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroB = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_signProd = mulAddRecFNToRaw_preMul_io_toPostMul_signProd; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isNaNC = mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isInfC = mulAddRecFNToRaw_preMul_io_toPostMul_isInfC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_isZeroC = mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_sExpSum = mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_doSubMags = mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CIsDominant = mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_CDom_CAlignDist = mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_highAlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_fromPreMul_bit0AlignedSigC = mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC; // @[MulAddRecFN.scala 332:44]
  assign mulAddRecFNToRaw_postMul_io_mulAddResult = _T + mulAddRecFNToRaw_preMul_io_mulAddC; // @[MulAddRecFN.scala 334:46]
  assign roundRawFNToRecFN_io_invalidExc = mulAddRecFNToRaw_postMul_io_invalidExc; // @[MulAddRecFN.scala 341:39]
  assign roundRawFNToRecFN_io_in_isNaN = mulAddRecFNToRaw_postMul_io_rawOut_isNaN; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isInf = mulAddRecFNToRaw_postMul_io_rawOut_isInf; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_isZero = mulAddRecFNToRaw_postMul_io_rawOut_isZero; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sign = mulAddRecFNToRaw_postMul_io_rawOut_sign; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sExp = mulAddRecFNToRaw_postMul_io_rawOut_sExp; // @[MulAddRecFN.scala 343:39]
  assign roundRawFNToRecFN_io_in_sig = mulAddRecFNToRaw_postMul_io_rawOut_sig; // @[MulAddRecFN.scala 343:39]
endmodule
module FPUALU(
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out
);
  wire [63:0] dummy1_io_in; // @[FPALU.scala 167:22]
  wire [64:0] dummy1_io_out; // @[FPALU.scala 167:22]
  wire [63:0] dummy0_io_in; // @[FPALU.scala 173:22]
  wire [64:0] dummy0_io_out; // @[FPALU.scala 173:22]
  wire [64:0] mulAddRecFN_io_a; // @[FPALU.scala 183:27]
  wire [64:0] mulAddRecFN_io_b; // @[FPALU.scala 183:27]
  wire [64:0] mulAddRecFN_io_c; // @[FPALU.scala 183:27]
  wire [64:0] mulAddRecFN_io_out; // @[FPALU.scala 183:27]
  wire  _T_3 = io_in1[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_in1[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_57 = io_in1[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  wire [5:0] _T_58 = io_in1[2] ? 6'h31 : _T_57; // @[Mux.scala 47:69]
  wire [5:0] _T_59 = io_in1[3] ? 6'h30 : _T_58; // @[Mux.scala 47:69]
  wire [5:0] _T_60 = io_in1[4] ? 6'h2f : _T_59; // @[Mux.scala 47:69]
  wire [5:0] _T_61 = io_in1[5] ? 6'h2e : _T_60; // @[Mux.scala 47:69]
  wire [5:0] _T_62 = io_in1[6] ? 6'h2d : _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_63 = io_in1[7] ? 6'h2c : _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_64 = io_in1[8] ? 6'h2b : _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_65 = io_in1[9] ? 6'h2a : _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_66 = io_in1[10] ? 6'h29 : _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_67 = io_in1[11] ? 6'h28 : _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_68 = io_in1[12] ? 6'h27 : _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_69 = io_in1[13] ? 6'h26 : _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_70 = io_in1[14] ? 6'h25 : _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_71 = io_in1[15] ? 6'h24 : _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_72 = io_in1[16] ? 6'h23 : _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_73 = io_in1[17] ? 6'h22 : _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_74 = io_in1[18] ? 6'h21 : _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_75 = io_in1[19] ? 6'h20 : _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_76 = io_in1[20] ? 6'h1f : _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_77 = io_in1[21] ? 6'h1e : _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_78 = io_in1[22] ? 6'h1d : _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_79 = io_in1[23] ? 6'h1c : _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_80 = io_in1[24] ? 6'h1b : _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_81 = io_in1[25] ? 6'h1a : _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_82 = io_in1[26] ? 6'h19 : _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_83 = io_in1[27] ? 6'h18 : _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_84 = io_in1[28] ? 6'h17 : _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_85 = io_in1[29] ? 6'h16 : _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_86 = io_in1[30] ? 6'h15 : _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_87 = io_in1[31] ? 6'h14 : _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_88 = io_in1[32] ? 6'h13 : _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_89 = io_in1[33] ? 6'h12 : _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_90 = io_in1[34] ? 6'h11 : _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_91 = io_in1[35] ? 6'h10 : _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_92 = io_in1[36] ? 6'hf : _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_93 = io_in1[37] ? 6'he : _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_94 = io_in1[38] ? 6'hd : _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_95 = io_in1[39] ? 6'hc : _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_96 = io_in1[40] ? 6'hb : _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_97 = io_in1[41] ? 6'ha : _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_98 = io_in1[42] ? 6'h9 : _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_99 = io_in1[43] ? 6'h8 : _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_100 = io_in1[44] ? 6'h7 : _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_101 = io_in1[45] ? 6'h6 : _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_102 = io_in1[46] ? 6'h5 : _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_103 = io_in1[47] ? 6'h4 : _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_104 = io_in1[48] ? 6'h3 : _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_105 = io_in1[49] ? 6'h2 : _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_106 = io_in1[50] ? 6'h1 : _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_107 = io_in1[51] ? 6'h0 : _T_106; // @[Mux.scala 47:69]
  wire [114:0] _GEN_0 = {{63'd0}, io_in1[51:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_108 = _GEN_0 << _T_107; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_110 = {_T_108[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_1 = {{6'd0}, _T_107}; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_111 = _GEN_1 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_112 = _T_3 ? _T_111 : {{1'd0}, io_in1[62:52]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_113 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_2 = {{9'd0}, _T_113}; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_114 = 11'h400 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_3 = {{1'd0}, _T_114}; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_116 = _T_112 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_117 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_119 = _T_116[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_121 = ~_T_4; // @[rawFloatFromFN.scala 66:36]
  wire  _T_122 = _T_119 & _T_121; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_125 = {1'b0,$signed(_T_116)}; // @[rawFloatFromFN.scala 70:48]
  wire  _T_126 = ~_T_117; // @[rawFloatFromFN.scala 72:29]
  wire [51:0] _T_127 = _T_3 ? _T_110 : io_in1[51:0]; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_129 = {1'h0,_T_126,_T_127}; // @[Cat.scala 29:58]
  wire [2:0] _T_131 = _T_117 ? 3'h0 : _T_125[11:9]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_122}; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_133 = _T_131 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_136 = {_T_125[8:0],_T_129[51:0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_137 = {io_in1[63],_T_133}; // @[Cat.scala 29:58]
  wire  _T_141 = io_in2[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_142 = io_in2[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_195 = io_in2[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  wire [5:0] _T_196 = io_in2[2] ? 6'h31 : _T_195; // @[Mux.scala 47:69]
  wire [5:0] _T_197 = io_in2[3] ? 6'h30 : _T_196; // @[Mux.scala 47:69]
  wire [5:0] _T_198 = io_in2[4] ? 6'h2f : _T_197; // @[Mux.scala 47:69]
  wire [5:0] _T_199 = io_in2[5] ? 6'h2e : _T_198; // @[Mux.scala 47:69]
  wire [5:0] _T_200 = io_in2[6] ? 6'h2d : _T_199; // @[Mux.scala 47:69]
  wire [5:0] _T_201 = io_in2[7] ? 6'h2c : _T_200; // @[Mux.scala 47:69]
  wire [5:0] _T_202 = io_in2[8] ? 6'h2b : _T_201; // @[Mux.scala 47:69]
  wire [5:0] _T_203 = io_in2[9] ? 6'h2a : _T_202; // @[Mux.scala 47:69]
  wire [5:0] _T_204 = io_in2[10] ? 6'h29 : _T_203; // @[Mux.scala 47:69]
  wire [5:0] _T_205 = io_in2[11] ? 6'h28 : _T_204; // @[Mux.scala 47:69]
  wire [5:0] _T_206 = io_in2[12] ? 6'h27 : _T_205; // @[Mux.scala 47:69]
  wire [5:0] _T_207 = io_in2[13] ? 6'h26 : _T_206; // @[Mux.scala 47:69]
  wire [5:0] _T_208 = io_in2[14] ? 6'h25 : _T_207; // @[Mux.scala 47:69]
  wire [5:0] _T_209 = io_in2[15] ? 6'h24 : _T_208; // @[Mux.scala 47:69]
  wire [5:0] _T_210 = io_in2[16] ? 6'h23 : _T_209; // @[Mux.scala 47:69]
  wire [5:0] _T_211 = io_in2[17] ? 6'h22 : _T_210; // @[Mux.scala 47:69]
  wire [5:0] _T_212 = io_in2[18] ? 6'h21 : _T_211; // @[Mux.scala 47:69]
  wire [5:0] _T_213 = io_in2[19] ? 6'h20 : _T_212; // @[Mux.scala 47:69]
  wire [5:0] _T_214 = io_in2[20] ? 6'h1f : _T_213; // @[Mux.scala 47:69]
  wire [5:0] _T_215 = io_in2[21] ? 6'h1e : _T_214; // @[Mux.scala 47:69]
  wire [5:0] _T_216 = io_in2[22] ? 6'h1d : _T_215; // @[Mux.scala 47:69]
  wire [5:0] _T_217 = io_in2[23] ? 6'h1c : _T_216; // @[Mux.scala 47:69]
  wire [5:0] _T_218 = io_in2[24] ? 6'h1b : _T_217; // @[Mux.scala 47:69]
  wire [5:0] _T_219 = io_in2[25] ? 6'h1a : _T_218; // @[Mux.scala 47:69]
  wire [5:0] _T_220 = io_in2[26] ? 6'h19 : _T_219; // @[Mux.scala 47:69]
  wire [5:0] _T_221 = io_in2[27] ? 6'h18 : _T_220; // @[Mux.scala 47:69]
  wire [5:0] _T_222 = io_in2[28] ? 6'h17 : _T_221; // @[Mux.scala 47:69]
  wire [5:0] _T_223 = io_in2[29] ? 6'h16 : _T_222; // @[Mux.scala 47:69]
  wire [5:0] _T_224 = io_in2[30] ? 6'h15 : _T_223; // @[Mux.scala 47:69]
  wire [5:0] _T_225 = io_in2[31] ? 6'h14 : _T_224; // @[Mux.scala 47:69]
  wire [5:0] _T_226 = io_in2[32] ? 6'h13 : _T_225; // @[Mux.scala 47:69]
  wire [5:0] _T_227 = io_in2[33] ? 6'h12 : _T_226; // @[Mux.scala 47:69]
  wire [5:0] _T_228 = io_in2[34] ? 6'h11 : _T_227; // @[Mux.scala 47:69]
  wire [5:0] _T_229 = io_in2[35] ? 6'h10 : _T_228; // @[Mux.scala 47:69]
  wire [5:0] _T_230 = io_in2[36] ? 6'hf : _T_229; // @[Mux.scala 47:69]
  wire [5:0] _T_231 = io_in2[37] ? 6'he : _T_230; // @[Mux.scala 47:69]
  wire [5:0] _T_232 = io_in2[38] ? 6'hd : _T_231; // @[Mux.scala 47:69]
  wire [5:0] _T_233 = io_in2[39] ? 6'hc : _T_232; // @[Mux.scala 47:69]
  wire [5:0] _T_234 = io_in2[40] ? 6'hb : _T_233; // @[Mux.scala 47:69]
  wire [5:0] _T_235 = io_in2[41] ? 6'ha : _T_234; // @[Mux.scala 47:69]
  wire [5:0] _T_236 = io_in2[42] ? 6'h9 : _T_235; // @[Mux.scala 47:69]
  wire [5:0] _T_237 = io_in2[43] ? 6'h8 : _T_236; // @[Mux.scala 47:69]
  wire [5:0] _T_238 = io_in2[44] ? 6'h7 : _T_237; // @[Mux.scala 47:69]
  wire [5:0] _T_239 = io_in2[45] ? 6'h6 : _T_238; // @[Mux.scala 47:69]
  wire [5:0] _T_240 = io_in2[46] ? 6'h5 : _T_239; // @[Mux.scala 47:69]
  wire [5:0] _T_241 = io_in2[47] ? 6'h4 : _T_240; // @[Mux.scala 47:69]
  wire [5:0] _T_242 = io_in2[48] ? 6'h3 : _T_241; // @[Mux.scala 47:69]
  wire [5:0] _T_243 = io_in2[49] ? 6'h2 : _T_242; // @[Mux.scala 47:69]
  wire [5:0] _T_244 = io_in2[50] ? 6'h1 : _T_243; // @[Mux.scala 47:69]
  wire [5:0] _T_245 = io_in2[51] ? 6'h0 : _T_244; // @[Mux.scala 47:69]
  wire [114:0] _GEN_5 = {{63'd0}, io_in2[51:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_246 = _GEN_5 << _T_245; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_248 = {_T_246[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_6 = {{6'd0}, _T_245}; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_249 = _GEN_6 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_250 = _T_141 ? _T_249 : {{1'd0}, io_in2[62:52]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_251 = _T_141 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_7 = {{9'd0}, _T_251}; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_252 = 11'h400 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_8 = {{1'd0}, _T_252}; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_254 = _T_250 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_255 = _T_141 & _T_142; // @[rawFloatFromFN.scala 62:34]
  wire  _T_257 = _T_254[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_259 = ~_T_142; // @[rawFloatFromFN.scala 66:36]
  wire  _T_260 = _T_257 & _T_259; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_263 = {1'b0,$signed(_T_254)}; // @[rawFloatFromFN.scala 70:48]
  wire  _T_264 = ~_T_255; // @[rawFloatFromFN.scala 72:29]
  wire [51:0] _T_265 = _T_141 ? _T_248 : io_in2[51:0]; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_267 = {1'h0,_T_264,_T_265}; // @[Cat.scala 29:58]
  wire [2:0] _T_269 = _T_255 ? 3'h0 : _T_263[11:9]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_260}; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_271 = _T_269 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_274 = {_T_263[8:0],_T_267[51:0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_275 = {io_in2[63],_T_271}; // @[Cat.scala 29:58]
  wire  _T_278 = mulAddRecFN_io_out[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_280 = mulAddRecFN_io_out[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_283 = _T_280 & mulAddRecFN_io_out[61]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_285 = ~mulAddRecFN_io_out[61]; // @[rawFloatFromRecFN.scala 56:36]
  wire  _T_286 = _T_280 & _T_285; // @[rawFloatFromRecFN.scala 56:33]
  wire [12:0] _T_288 = {1'b0,$signed(mulAddRecFN_io_out[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _T_289 = ~_T_278; // @[rawFloatFromRecFN.scala 60:39]
  wire [53:0] _T_292 = {1'h0,_T_289,mulAddRecFN_io_out[51:0]}; // @[Cat.scala 29:58]
  wire  _T_293 = $signed(_T_288) < 13'sh402; // @[fNFromRecFN.scala 50:39]
  wire [5:0] _T_296 = 6'h1 - _T_288[5:0]; // @[fNFromRecFN.scala 51:39]
  wire [52:0] _T_298 = _T_292[53:1] >> _T_296; // @[fNFromRecFN.scala 52:42]
  wire [10:0] _T_302 = _T_288[10:0] - 11'h401; // @[fNFromRecFN.scala 57:45]
  wire [10:0] _T_303 = _T_293 ? 11'h0 : _T_302; // @[fNFromRecFN.scala 55:16]
  wire  _T_304 = _T_283 | _T_286; // @[fNFromRecFN.scala 59:44]
  wire [10:0] _T_306 = _T_304 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _T_307 = _T_303 | _T_306; // @[fNFromRecFN.scala 59:15]
  wire [51:0] _T_309 = _T_286 ? 52'h0 : _T_292[51:0]; // @[fNFromRecFN.scala 63:20]
  wire [51:0] _T_310 = _T_293 ? _T_298[51:0] : _T_309; // @[fNFromRecFN.scala 61:16]
  wire [11:0] _T_311 = {mulAddRecFN_io_out[64],_T_307}; // @[Cat.scala 29:58]
  INToRecFN dummy1 ( // @[FPALU.scala 167:22]
    .io_in(dummy1_io_in),
    .io_out(dummy1_io_out)
  );
  INToRecFN dummy0 ( // @[FPALU.scala 173:22]
    .io_in(dummy0_io_in),
    .io_out(dummy0_io_out)
  );
  MulAddRecFN mulAddRecFN ( // @[FPALU.scala 183:27]
    .io_a(mulAddRecFN_io_a),
    .io_b(mulAddRecFN_io_b),
    .io_c(mulAddRecFN_io_c),
    .io_out(mulAddRecFN_io_out)
  );
  assign io_out = {_T_311,_T_310}; // @[FPALU.scala 190:10]
  assign dummy1_io_in = 64'h1; // @[FPALU.scala 169:16]
  assign dummy0_io_in = 64'h0; // @[FPALU.scala 175:16]
  assign mulAddRecFN_io_a = {_T_137,_T_136}; // @[FPALU.scala 150:26]
  assign mulAddRecFN_io_b = {_T_275,_T_274}; // @[FPALU.scala 151:26]
  assign mulAddRecFN_io_c = dummy0_io_out; // @[FPALU.scala 152:26]
endmodule
module FPComputeNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[FPComputeNode.scala 64:18]
  wire [63:0] FU_io_in2; // @[FPComputeNode.scala 64:18]
  wire [63:0] FU_io_out; // @[FPComputeNode.scala 64:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [63:0] left_R_data; // @[FPComputeNode.scala 51:23]
  reg  left_valid_R; // @[FPComputeNode.scala 52:29]
  reg [63:0] right_R_data; // @[FPComputeNode.scala 55:24]
  reg  right_valid_R; // @[FPComputeNode.scala 56:30]
  reg [4:0] task_ID_R; // @[FPComputeNode.scala 58:26]
  reg  state; // @[FPComputeNode.scala 62:22]
  reg [63:0] out_data_R; // @[FPComputeNode.scala 66:27]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[FPComputeNode.scala 79:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[FPComputeNode.scala 85:27]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & left_valid_R; // @[FPComputeNode.scala 99:27]
  wire  _T_18 = _T_17 & right_valid_R; // @[FPComputeNode.scala 99:43]
  wire  _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire [14:0] _T_24 = value + 15'h1; // @[Counter.scala 39:22]
  wire  _T_26 = ~reset; // @[FPComputeNode.scala 108:17]
  wire [63:0] _T_19_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_16 = _T_18 ? _T_19_data : out_data_R; // @[FPComputeNode.scala 99:61]
  wire  _GEN_19 = _T_18 | out_valid_R_0; // @[FPComputeNode.scala 99:61]
  wire  _GEN_23 = _T_18 | state; // @[FPComputeNode.scala 99:61]
  wire  _T_29 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_45 = _T_16 & _T_18; // @[FPComputeNode.scala 108:17]
  FPUALU FU ( // @[FPComputeNode.scala 64:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_16 ? _GEN_19 : out_valid_R_0; // @[HandShaking.scala 194:21 FPComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_16 : out_data_R; // @[FPComputeNode.scala 92:25 FPComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~left_valid_R; // @[FPComputeNode.scala 78:19]
  assign io_RightIO_ready = ~right_valid_R; // @[FPComputeNode.scala 84:20]
  assign FU_io_in1 = left_R_data; // @[FPComputeNode.scala 75:13]
  assign FU_io_in2 = right_R_data; // @[FPComputeNode.scala 76:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[14:0];
  _RAND_7 = {2{`RANDOM}};
  left_R_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  left_valid_R = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  right_R_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  task_ID_R = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_29) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_16) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_29) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        out_valid_R_0 <= _T_21;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      value <= 15'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        value <= _T_24;
      end
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    task_ID_R <= enable_R_taskID;
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_23;
    end else if (state) begin
      if (_T_29) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_16) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_29) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_45 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [FPCompute] [FP_mul2121] [Pred: %d] [Iter: %d] [In(0): %d] [In(1) %d] [Out: %d] [OpCode: fmul] [Cycle: %d]\n",task_ID_R,enable_R_control,value,left_R_data,right_R_data,FU_io_out,cycleCount); // @[FPComputeNode.scala 108:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_22] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_23] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [63:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [63:0] io_idx_0_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_ready_R_1; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  reg  out_valid_R_1; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_8 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] base_addr_R_data; // @[GepNode.scala 884:28]
  reg  base_addr_valid_R; // @[GepNode.scala 885:34]
  reg [63:0] idx_R_0_data; // @[GepNode.scala 888:39]
  reg  idx_valid_R_0; // @[GepNode.scala 889:45]
  reg  state; // @[GepNode.scala 893:22]
  wire  _T_12 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_12 | base_addr_valid_R; // @[GepNode.scala 909:31]
  wire  _T_14 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_14 | idx_valid_R_0; // @[GepNode.scala 916:28]
  wire [67:0] seek_value = idx_R_0_data * 64'h8; // @[GepNode.scala 924:21]
  wire [67:0] _GEN_59 = {{4'd0}, base_addr_R_data}; // @[GepNode.scala 932:35]
  wire [67:0] data_out = _GEN_59 + seek_value; // @[GepNode.scala 932:35]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 948:27]
  wire  _T_18 = _T_17 & idx_valid_R_0; // @[GepNode.scala 948:48]
  wire  _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_22 = _T_2 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _GEN_20 = _T_18 | state; // @[GepNode.scala 948:78]
  wire  _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_27 = out_ready_R_1 | _T_2; // @[HandShaking.scala 251:83]
  wire  _T_28 = _T_26 & _T_27; // @[HandShaking.scala 252:27]
  wire  _T_32 = ~reset; // @[GepNode.scala 968:17]
  wire  _GEN_60 = ~_T_16; // @[GepNode.scala 968:17]
  wire  _GEN_61 = _GEN_60 & state; // @[GepNode.scala 968:17]
  wire  _GEN_62 = _GEN_61 & _T_28; // @[GepNode.scala 968:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 194:21]
  assign io_Out_0_bits_data = data_out[63:0]; // @[GepNode.scala 936:25]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 194:21]
  assign io_Out_1_bits_data = data_out[63:0]; // @[GepNode.scala 936:25]
  assign io_baseAddress_ready = ~base_addr_valid_R; // @[GepNode.scala 908:24]
  assign io_idx_0_ready = ~idx_valid_R_0; // @[GepNode.scala 915:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {2{`RANDOM}};
  base_addr_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  idx_R_0_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_4) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_4) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_28) begin
        enable_valid_R <= 1'h0;
      end else if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_4) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_16) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_28) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_16) begin
      if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_28) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_2) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        out_valid_R_0 <= _T_21;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        out_valid_R_1 <= _T_22;
      end else if (_T_2) begin
        out_valid_R_1 <= 1'h0;
      end
    end else if (_T_2) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_8;
    end
    if (reset) begin
      base_addr_R_data <= 64'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        base_addr_R_data <= io_baseAddress_bits_data;
      end
    end else if (state) begin
      if (_T_28) begin
        base_addr_R_data <= 64'h0;
      end else if (_T_12) begin
        base_addr_R_data <= io_baseAddress_bits_data;
      end
    end else if (_T_12) begin
      base_addr_R_data <= io_baseAddress_bits_data;
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else if (_T_16) begin
      base_addr_valid_R <= _GEN_13;
    end else if (state) begin
      if (_T_28) begin
        base_addr_valid_R <= 1'h0;
      end else begin
        base_addr_valid_R <= _GEN_13;
      end
    end else begin
      base_addr_valid_R <= _GEN_13;
    end
    if (reset) begin
      idx_R_0_data <= 64'h0;
    end else if (_T_16) begin
      if (_T_14) begin
        idx_R_0_data <= io_idx_0_bits_data;
      end
    end else if (state) begin
      if (_T_28) begin
        idx_R_0_data <= 64'h0;
      end else if (_T_14) begin
        idx_R_0_data <= io_idx_0_bits_data;
      end
    end else if (_T_14) begin
      idx_R_0_data <= io_idx_0_bits_data;
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      idx_valid_R_0 <= _GEN_17;
    end else if (state) begin
      if (_T_28) begin
        idx_valid_R_0 <= 1'h0;
      end else begin
        idx_valid_R_0 <= _GEN_17;
      end
    end else begin
      idx_valid_R_0 <= _GEN_17;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_20;
    end else if (state) begin
      if (_T_28) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_32) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [GEP] [Gep_arrayidx2524] [Pred: %d][Out: 0x%x] [Cycle: %d]\n",enable_R_taskID,enable_R_control,data_out,cycleCount); // @[GepNode.scala 968:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoadCache_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [63:0] io_GepAddr_bits_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [63:0] io_MemReq_bits_addr,
  input         io_MemResp_valid,
  input  [63:0] io_MemResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  out_ready_R_0; // @[HandShaking.scala 605:28]
  reg  out_valid_R_0; // @[HandShaking.scala 606:28]
  wire  _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_4 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 632:29]
  wire  _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_10 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [63:0] addr_R_data; // @[LoadCache.scala 58:23]
  reg  addr_valid_R; // @[LoadCache.scala 59:29]
  reg [63:0] data_R_data; // @[LoadCache.scala 62:23]
  reg [1:0] state; // @[LoadCache.scala 67:22]
  wire  _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_14 | addr_valid_R; // @[LoadCache.scala 76:27]
  wire  _T_15 = enable_valid_R & addr_valid_R; // @[LoadCache.scala 95:20]
  wire  _T_16 = _T_15 & enable_R_control; // @[LoadCache.scala 95:36]
  wire  _T_23 = &out_ready_R_0; // @[HandShaking.scala 725:24]
  wire  _T_24 = &io_Out_0_ready; // @[HandShaking.scala 725:50]
  wire  _T_25 = _T_23 | _T_24; // @[HandShaking.scala 725:29]
  wire  _T_44 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_49 = _T_4 ^ 1'h1; // @[HandShaking.scala 729:72]
  wire  _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_25 = io_MemResp_valid | _GEN_1; // @[LoadCache.scala 214:30]
  wire  _T_51 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [14:0] _T_62 = value + 15'h1; // @[Counter.scala 39:22]
  wire  _T_64 = ~reset; // @[LoadCache.scala 254:17]
  wire  _GEN_78 = ~_T_44; // @[LoadCache.scala 254:17]
  wire  _GEN_79 = ~_T_50; // @[LoadCache.scala 254:17]
  wire  _GEN_80 = _GEN_78 & _GEN_79; // @[LoadCache.scala 254:17]
  wire  _GEN_81 = _GEN_80 & _T_51; // @[LoadCache.scala 254:17]
  wire  _GEN_82 = _GEN_81 & _T_25; // @[LoadCache.scala 254:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 630:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadCache.scala 158:20]
  assign io_GepAddr_ready = ~addr_valid_R; // @[LoadCache.scala 75:20]
  assign io_MemReq_valid = _T_44 & _T_16; // @[LoadCache.scala 162:19 LoadCache.scala 185:27]
  assign io_MemReq_bits_addr = addr_R_data; // @[LoadCache.scala 164:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[14:0];
  _RAND_7 = {2{`RANDOM}};
  addr_R_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  data_R_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_6) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_6) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_44) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_50) begin
      if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_44) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_50) begin
      if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_4) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_4) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_44) begin
      if (_T_15) begin
        if (enable_R_control) begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end else begin
          out_valid_R_0 <= _T_49;
        end
      end else if (_T_4) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_50) begin
      out_valid_R_0 <= _GEN_25;
    end else if (_T_4) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_10;
    end
    if (reset) begin
      value <= 15'h0;
    end else if (!(_T_44)) begin
      if (!(_T_50)) begin
        if (_T_51) begin
          if (_T_25) begin
            value <= _T_62;
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 64'h0;
    end else if (_T_44) begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_50) begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        addr_R_data <= 64'h0;
      end else if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_14) begin
      addr_R_data <= io_GepAddr_bits_data;
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else if (_T_44) begin
      addr_valid_R <= _GEN_11;
    end else if (_T_50) begin
      addr_valid_R <= _GEN_11;
    end else if (_T_51) begin
      if (_T_25) begin
        addr_valid_R <= 1'h0;
      end else begin
        addr_valid_R <= _GEN_11;
      end
    end else begin
      addr_valid_R <= _GEN_11;
    end
    if (reset) begin
      data_R_data <= 64'h0;
    end else if (!(_T_44)) begin
      if (_T_50) begin
        if (io_MemResp_valid) begin
          data_R_data <= io_MemResp_bits_data;
        end
      end else if (_T_51) begin
        if (_T_25) begin
          data_R_data <= 64'h0;
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_44) begin
      if (_T_15) begin
        if (enable_R_control) begin
          if (io_MemReq_ready) begin
            state <= 2'h1;
          end
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_50) begin
      if (io_MemResp_valid) begin
        state <= 2'h2;
      end
    end else if (_T_51) begin
      if (_T_25) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [LOAD] [ld_25] [Pred: %d] [Iter: %d] [Addr: %d] [Data: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,value,addr_R_data,data_R_data,cycleCount); // @[LoadCache.scala 254:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module FPUALU_1(
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out
);
  wire [63:0] dummy1_io_in; // @[FPALU.scala 167:22]
  wire [64:0] dummy1_io_out; // @[FPALU.scala 167:22]
  wire [63:0] dummy0_io_in; // @[FPALU.scala 173:22]
  wire [64:0] dummy0_io_out; // @[FPALU.scala 173:22]
  wire [64:0] mulAddRecFN_io_a; // @[FPALU.scala 183:27]
  wire [64:0] mulAddRecFN_io_b; // @[FPALU.scala 183:27]
  wire [64:0] mulAddRecFN_io_c; // @[FPALU.scala 183:27]
  wire [64:0] mulAddRecFN_io_out; // @[FPALU.scala 183:27]
  wire  _T_3 = io_in1[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_4 = io_in1[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_57 = io_in1[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  wire [5:0] _T_58 = io_in1[2] ? 6'h31 : _T_57; // @[Mux.scala 47:69]
  wire [5:0] _T_59 = io_in1[3] ? 6'h30 : _T_58; // @[Mux.scala 47:69]
  wire [5:0] _T_60 = io_in1[4] ? 6'h2f : _T_59; // @[Mux.scala 47:69]
  wire [5:0] _T_61 = io_in1[5] ? 6'h2e : _T_60; // @[Mux.scala 47:69]
  wire [5:0] _T_62 = io_in1[6] ? 6'h2d : _T_61; // @[Mux.scala 47:69]
  wire [5:0] _T_63 = io_in1[7] ? 6'h2c : _T_62; // @[Mux.scala 47:69]
  wire [5:0] _T_64 = io_in1[8] ? 6'h2b : _T_63; // @[Mux.scala 47:69]
  wire [5:0] _T_65 = io_in1[9] ? 6'h2a : _T_64; // @[Mux.scala 47:69]
  wire [5:0] _T_66 = io_in1[10] ? 6'h29 : _T_65; // @[Mux.scala 47:69]
  wire [5:0] _T_67 = io_in1[11] ? 6'h28 : _T_66; // @[Mux.scala 47:69]
  wire [5:0] _T_68 = io_in1[12] ? 6'h27 : _T_67; // @[Mux.scala 47:69]
  wire [5:0] _T_69 = io_in1[13] ? 6'h26 : _T_68; // @[Mux.scala 47:69]
  wire [5:0] _T_70 = io_in1[14] ? 6'h25 : _T_69; // @[Mux.scala 47:69]
  wire [5:0] _T_71 = io_in1[15] ? 6'h24 : _T_70; // @[Mux.scala 47:69]
  wire [5:0] _T_72 = io_in1[16] ? 6'h23 : _T_71; // @[Mux.scala 47:69]
  wire [5:0] _T_73 = io_in1[17] ? 6'h22 : _T_72; // @[Mux.scala 47:69]
  wire [5:0] _T_74 = io_in1[18] ? 6'h21 : _T_73; // @[Mux.scala 47:69]
  wire [5:0] _T_75 = io_in1[19] ? 6'h20 : _T_74; // @[Mux.scala 47:69]
  wire [5:0] _T_76 = io_in1[20] ? 6'h1f : _T_75; // @[Mux.scala 47:69]
  wire [5:0] _T_77 = io_in1[21] ? 6'h1e : _T_76; // @[Mux.scala 47:69]
  wire [5:0] _T_78 = io_in1[22] ? 6'h1d : _T_77; // @[Mux.scala 47:69]
  wire [5:0] _T_79 = io_in1[23] ? 6'h1c : _T_78; // @[Mux.scala 47:69]
  wire [5:0] _T_80 = io_in1[24] ? 6'h1b : _T_79; // @[Mux.scala 47:69]
  wire [5:0] _T_81 = io_in1[25] ? 6'h1a : _T_80; // @[Mux.scala 47:69]
  wire [5:0] _T_82 = io_in1[26] ? 6'h19 : _T_81; // @[Mux.scala 47:69]
  wire [5:0] _T_83 = io_in1[27] ? 6'h18 : _T_82; // @[Mux.scala 47:69]
  wire [5:0] _T_84 = io_in1[28] ? 6'h17 : _T_83; // @[Mux.scala 47:69]
  wire [5:0] _T_85 = io_in1[29] ? 6'h16 : _T_84; // @[Mux.scala 47:69]
  wire [5:0] _T_86 = io_in1[30] ? 6'h15 : _T_85; // @[Mux.scala 47:69]
  wire [5:0] _T_87 = io_in1[31] ? 6'h14 : _T_86; // @[Mux.scala 47:69]
  wire [5:0] _T_88 = io_in1[32] ? 6'h13 : _T_87; // @[Mux.scala 47:69]
  wire [5:0] _T_89 = io_in1[33] ? 6'h12 : _T_88; // @[Mux.scala 47:69]
  wire [5:0] _T_90 = io_in1[34] ? 6'h11 : _T_89; // @[Mux.scala 47:69]
  wire [5:0] _T_91 = io_in1[35] ? 6'h10 : _T_90; // @[Mux.scala 47:69]
  wire [5:0] _T_92 = io_in1[36] ? 6'hf : _T_91; // @[Mux.scala 47:69]
  wire [5:0] _T_93 = io_in1[37] ? 6'he : _T_92; // @[Mux.scala 47:69]
  wire [5:0] _T_94 = io_in1[38] ? 6'hd : _T_93; // @[Mux.scala 47:69]
  wire [5:0] _T_95 = io_in1[39] ? 6'hc : _T_94; // @[Mux.scala 47:69]
  wire [5:0] _T_96 = io_in1[40] ? 6'hb : _T_95; // @[Mux.scala 47:69]
  wire [5:0] _T_97 = io_in1[41] ? 6'ha : _T_96; // @[Mux.scala 47:69]
  wire [5:0] _T_98 = io_in1[42] ? 6'h9 : _T_97; // @[Mux.scala 47:69]
  wire [5:0] _T_99 = io_in1[43] ? 6'h8 : _T_98; // @[Mux.scala 47:69]
  wire [5:0] _T_100 = io_in1[44] ? 6'h7 : _T_99; // @[Mux.scala 47:69]
  wire [5:0] _T_101 = io_in1[45] ? 6'h6 : _T_100; // @[Mux.scala 47:69]
  wire [5:0] _T_102 = io_in1[46] ? 6'h5 : _T_101; // @[Mux.scala 47:69]
  wire [5:0] _T_103 = io_in1[47] ? 6'h4 : _T_102; // @[Mux.scala 47:69]
  wire [5:0] _T_104 = io_in1[48] ? 6'h3 : _T_103; // @[Mux.scala 47:69]
  wire [5:0] _T_105 = io_in1[49] ? 6'h2 : _T_104; // @[Mux.scala 47:69]
  wire [5:0] _T_106 = io_in1[50] ? 6'h1 : _T_105; // @[Mux.scala 47:69]
  wire [5:0] _T_107 = io_in1[51] ? 6'h0 : _T_106; // @[Mux.scala 47:69]
  wire [114:0] _GEN_0 = {{63'd0}, io_in1[51:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_108 = _GEN_0 << _T_107; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_110 = {_T_108[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_1 = {{6'd0}, _T_107}; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_111 = _GEN_1 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_112 = _T_3 ? _T_111 : {{1'd0}, io_in1[62:52]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_113 = _T_3 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_2 = {{9'd0}, _T_113}; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_114 = 11'h400 | _GEN_2; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_3 = {{1'd0}, _T_114}; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_116 = _T_112 + _GEN_3; // @[rawFloatFromFN.scala 59:15]
  wire  _T_117 = _T_3 & _T_4; // @[rawFloatFromFN.scala 62:34]
  wire  _T_119 = _T_116[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_121 = ~_T_4; // @[rawFloatFromFN.scala 66:36]
  wire  _T_122 = _T_119 & _T_121; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_125 = {1'b0,$signed(_T_116)}; // @[rawFloatFromFN.scala 70:48]
  wire  _T_126 = ~_T_117; // @[rawFloatFromFN.scala 72:29]
  wire [51:0] _T_127 = _T_3 ? _T_110 : io_in1[51:0]; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_129 = {1'h0,_T_126,_T_127}; // @[Cat.scala 29:58]
  wire [2:0] _T_131 = _T_117 ? 3'h0 : _T_125[11:9]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_4 = {{2'd0}, _T_122}; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_133 = _T_131 | _GEN_4; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_136 = {_T_125[8:0],_T_129[51:0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_137 = {io_in1[63],_T_133}; // @[Cat.scala 29:58]
  wire  _T_141 = io_in2[62:52] == 11'h0; // @[rawFloatFromFN.scala 50:34]
  wire  _T_142 = io_in2[51:0] == 52'h0; // @[rawFloatFromFN.scala 51:38]
  wire [5:0] _T_195 = io_in2[1] ? 6'h32 : 6'h33; // @[Mux.scala 47:69]
  wire [5:0] _T_196 = io_in2[2] ? 6'h31 : _T_195; // @[Mux.scala 47:69]
  wire [5:0] _T_197 = io_in2[3] ? 6'h30 : _T_196; // @[Mux.scala 47:69]
  wire [5:0] _T_198 = io_in2[4] ? 6'h2f : _T_197; // @[Mux.scala 47:69]
  wire [5:0] _T_199 = io_in2[5] ? 6'h2e : _T_198; // @[Mux.scala 47:69]
  wire [5:0] _T_200 = io_in2[6] ? 6'h2d : _T_199; // @[Mux.scala 47:69]
  wire [5:0] _T_201 = io_in2[7] ? 6'h2c : _T_200; // @[Mux.scala 47:69]
  wire [5:0] _T_202 = io_in2[8] ? 6'h2b : _T_201; // @[Mux.scala 47:69]
  wire [5:0] _T_203 = io_in2[9] ? 6'h2a : _T_202; // @[Mux.scala 47:69]
  wire [5:0] _T_204 = io_in2[10] ? 6'h29 : _T_203; // @[Mux.scala 47:69]
  wire [5:0] _T_205 = io_in2[11] ? 6'h28 : _T_204; // @[Mux.scala 47:69]
  wire [5:0] _T_206 = io_in2[12] ? 6'h27 : _T_205; // @[Mux.scala 47:69]
  wire [5:0] _T_207 = io_in2[13] ? 6'h26 : _T_206; // @[Mux.scala 47:69]
  wire [5:0] _T_208 = io_in2[14] ? 6'h25 : _T_207; // @[Mux.scala 47:69]
  wire [5:0] _T_209 = io_in2[15] ? 6'h24 : _T_208; // @[Mux.scala 47:69]
  wire [5:0] _T_210 = io_in2[16] ? 6'h23 : _T_209; // @[Mux.scala 47:69]
  wire [5:0] _T_211 = io_in2[17] ? 6'h22 : _T_210; // @[Mux.scala 47:69]
  wire [5:0] _T_212 = io_in2[18] ? 6'h21 : _T_211; // @[Mux.scala 47:69]
  wire [5:0] _T_213 = io_in2[19] ? 6'h20 : _T_212; // @[Mux.scala 47:69]
  wire [5:0] _T_214 = io_in2[20] ? 6'h1f : _T_213; // @[Mux.scala 47:69]
  wire [5:0] _T_215 = io_in2[21] ? 6'h1e : _T_214; // @[Mux.scala 47:69]
  wire [5:0] _T_216 = io_in2[22] ? 6'h1d : _T_215; // @[Mux.scala 47:69]
  wire [5:0] _T_217 = io_in2[23] ? 6'h1c : _T_216; // @[Mux.scala 47:69]
  wire [5:0] _T_218 = io_in2[24] ? 6'h1b : _T_217; // @[Mux.scala 47:69]
  wire [5:0] _T_219 = io_in2[25] ? 6'h1a : _T_218; // @[Mux.scala 47:69]
  wire [5:0] _T_220 = io_in2[26] ? 6'h19 : _T_219; // @[Mux.scala 47:69]
  wire [5:0] _T_221 = io_in2[27] ? 6'h18 : _T_220; // @[Mux.scala 47:69]
  wire [5:0] _T_222 = io_in2[28] ? 6'h17 : _T_221; // @[Mux.scala 47:69]
  wire [5:0] _T_223 = io_in2[29] ? 6'h16 : _T_222; // @[Mux.scala 47:69]
  wire [5:0] _T_224 = io_in2[30] ? 6'h15 : _T_223; // @[Mux.scala 47:69]
  wire [5:0] _T_225 = io_in2[31] ? 6'h14 : _T_224; // @[Mux.scala 47:69]
  wire [5:0] _T_226 = io_in2[32] ? 6'h13 : _T_225; // @[Mux.scala 47:69]
  wire [5:0] _T_227 = io_in2[33] ? 6'h12 : _T_226; // @[Mux.scala 47:69]
  wire [5:0] _T_228 = io_in2[34] ? 6'h11 : _T_227; // @[Mux.scala 47:69]
  wire [5:0] _T_229 = io_in2[35] ? 6'h10 : _T_228; // @[Mux.scala 47:69]
  wire [5:0] _T_230 = io_in2[36] ? 6'hf : _T_229; // @[Mux.scala 47:69]
  wire [5:0] _T_231 = io_in2[37] ? 6'he : _T_230; // @[Mux.scala 47:69]
  wire [5:0] _T_232 = io_in2[38] ? 6'hd : _T_231; // @[Mux.scala 47:69]
  wire [5:0] _T_233 = io_in2[39] ? 6'hc : _T_232; // @[Mux.scala 47:69]
  wire [5:0] _T_234 = io_in2[40] ? 6'hb : _T_233; // @[Mux.scala 47:69]
  wire [5:0] _T_235 = io_in2[41] ? 6'ha : _T_234; // @[Mux.scala 47:69]
  wire [5:0] _T_236 = io_in2[42] ? 6'h9 : _T_235; // @[Mux.scala 47:69]
  wire [5:0] _T_237 = io_in2[43] ? 6'h8 : _T_236; // @[Mux.scala 47:69]
  wire [5:0] _T_238 = io_in2[44] ? 6'h7 : _T_237; // @[Mux.scala 47:69]
  wire [5:0] _T_239 = io_in2[45] ? 6'h6 : _T_238; // @[Mux.scala 47:69]
  wire [5:0] _T_240 = io_in2[46] ? 6'h5 : _T_239; // @[Mux.scala 47:69]
  wire [5:0] _T_241 = io_in2[47] ? 6'h4 : _T_240; // @[Mux.scala 47:69]
  wire [5:0] _T_242 = io_in2[48] ? 6'h3 : _T_241; // @[Mux.scala 47:69]
  wire [5:0] _T_243 = io_in2[49] ? 6'h2 : _T_242; // @[Mux.scala 47:69]
  wire [5:0] _T_244 = io_in2[50] ? 6'h1 : _T_243; // @[Mux.scala 47:69]
  wire [5:0] _T_245 = io_in2[51] ? 6'h0 : _T_244; // @[Mux.scala 47:69]
  wire [114:0] _GEN_5 = {{63'd0}, io_in2[51:0]}; // @[rawFloatFromFN.scala 54:36]
  wire [114:0] _T_246 = _GEN_5 << _T_245; // @[rawFloatFromFN.scala 54:36]
  wire [51:0] _T_248 = {_T_246[50:0], 1'h0}; // @[rawFloatFromFN.scala 54:64]
  wire [11:0] _GEN_6 = {{6'd0}, _T_245}; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_249 = _GEN_6 ^ 12'hfff; // @[rawFloatFromFN.scala 57:26]
  wire [11:0] _T_250 = _T_141 ? _T_249 : {{1'd0}, io_in2[62:52]}; // @[rawFloatFromFN.scala 56:16]
  wire [1:0] _T_251 = _T_141 ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 60:27]
  wire [10:0] _GEN_7 = {{9'd0}, _T_251}; // @[rawFloatFromFN.scala 60:22]
  wire [10:0] _T_252 = 11'h400 | _GEN_7; // @[rawFloatFromFN.scala 60:22]
  wire [11:0] _GEN_8 = {{1'd0}, _T_252}; // @[rawFloatFromFN.scala 59:15]
  wire [11:0] _T_254 = _T_250 + _GEN_8; // @[rawFloatFromFN.scala 59:15]
  wire  _T_255 = _T_141 & _T_142; // @[rawFloatFromFN.scala 62:34]
  wire  _T_257 = _T_254[11:10] == 2'h3; // @[rawFloatFromFN.scala 63:62]
  wire  _T_259 = ~_T_142; // @[rawFloatFromFN.scala 66:36]
  wire  _T_260 = _T_257 & _T_259; // @[rawFloatFromFN.scala 66:33]
  wire [12:0] _T_263 = {1'b0,$signed(_T_254)}; // @[rawFloatFromFN.scala 70:48]
  wire  _T_264 = ~_T_255; // @[rawFloatFromFN.scala 72:29]
  wire [51:0] _T_265 = _T_141 ? _T_248 : io_in2[51:0]; // @[rawFloatFromFN.scala 72:42]
  wire [53:0] _T_267 = {1'h0,_T_264,_T_265}; // @[Cat.scala 29:58]
  wire [2:0] _T_269 = _T_255 ? 3'h0 : _T_263[11:9]; // @[recFNFromFN.scala 48:16]
  wire [2:0] _GEN_9 = {{2'd0}, _T_260}; // @[recFNFromFN.scala 48:79]
  wire [2:0] _T_271 = _T_269 | _GEN_9; // @[recFNFromFN.scala 48:79]
  wire [60:0] _T_274 = {_T_263[8:0],_T_267[51:0]}; // @[Cat.scala 29:58]
  wire [3:0] _T_275 = {io_in2[63],_T_271}; // @[Cat.scala 29:58]
  wire  _T_278 = mulAddRecFN_io_out[63:61] == 3'h0; // @[rawFloatFromRecFN.scala 51:54]
  wire  _T_280 = mulAddRecFN_io_out[63:62] == 2'h3; // @[rawFloatFromRecFN.scala 52:54]
  wire  _T_283 = _T_280 & mulAddRecFN_io_out[61]; // @[rawFloatFromRecFN.scala 55:33]
  wire  _T_285 = ~mulAddRecFN_io_out[61]; // @[rawFloatFromRecFN.scala 56:36]
  wire  _T_286 = _T_280 & _T_285; // @[rawFloatFromRecFN.scala 56:33]
  wire [12:0] _T_288 = {1'b0,$signed(mulAddRecFN_io_out[63:52])}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _T_289 = ~_T_278; // @[rawFloatFromRecFN.scala 60:39]
  wire [53:0] _T_292 = {1'h0,_T_289,mulAddRecFN_io_out[51:0]}; // @[Cat.scala 29:58]
  wire  _T_293 = $signed(_T_288) < 13'sh402; // @[fNFromRecFN.scala 50:39]
  wire [5:0] _T_296 = 6'h1 - _T_288[5:0]; // @[fNFromRecFN.scala 51:39]
  wire [52:0] _T_298 = _T_292[53:1] >> _T_296; // @[fNFromRecFN.scala 52:42]
  wire [10:0] _T_302 = _T_288[10:0] - 11'h401; // @[fNFromRecFN.scala 57:45]
  wire [10:0] _T_303 = _T_293 ? 11'h0 : _T_302; // @[fNFromRecFN.scala 55:16]
  wire  _T_304 = _T_283 | _T_286; // @[fNFromRecFN.scala 59:44]
  wire [10:0] _T_306 = _T_304 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [10:0] _T_307 = _T_303 | _T_306; // @[fNFromRecFN.scala 59:15]
  wire [51:0] _T_309 = _T_286 ? 52'h0 : _T_292[51:0]; // @[fNFromRecFN.scala 63:20]
  wire [51:0] _T_310 = _T_293 ? _T_298[51:0] : _T_309; // @[fNFromRecFN.scala 61:16]
  wire [11:0] _T_311 = {mulAddRecFN_io_out[64],_T_307}; // @[Cat.scala 29:58]
  INToRecFN dummy1 ( // @[FPALU.scala 167:22]
    .io_in(dummy1_io_in),
    .io_out(dummy1_io_out)
  );
  INToRecFN dummy0 ( // @[FPALU.scala 173:22]
    .io_in(dummy0_io_in),
    .io_out(dummy0_io_out)
  );
  MulAddRecFN mulAddRecFN ( // @[FPALU.scala 183:27]
    .io_a(mulAddRecFN_io_a),
    .io_b(mulAddRecFN_io_b),
    .io_c(mulAddRecFN_io_c),
    .io_out(mulAddRecFN_io_out)
  );
  assign io_out = {_T_311,_T_310}; // @[FPALU.scala 190:10]
  assign dummy1_io_in = 64'h1; // @[FPALU.scala 169:16]
  assign dummy0_io_in = 64'h0; // @[FPALU.scala 175:16]
  assign mulAddRecFN_io_a = dummy1_io_out; // @[FPALU.scala 138:26]
  assign mulAddRecFN_io_b = {_T_137,_T_136}; // @[FPALU.scala 139:26]
  assign mulAddRecFN_io_c = {_T_275,_T_274}; // @[FPALU.scala 140:26]
endmodule
module FPComputeNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [63:0] io_RightIO_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[FPComputeNode.scala 64:18]
  wire [63:0] FU_io_in2; // @[FPComputeNode.scala 64:18]
  wire [63:0] FU_io_out; // @[FPComputeNode.scala 64:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [63:0] left_R_data; // @[FPComputeNode.scala 51:23]
  reg  left_valid_R; // @[FPComputeNode.scala 52:29]
  reg [63:0] right_R_data; // @[FPComputeNode.scala 55:24]
  reg  right_valid_R; // @[FPComputeNode.scala 56:30]
  reg [4:0] task_ID_R; // @[FPComputeNode.scala 58:26]
  reg  state; // @[FPComputeNode.scala 62:22]
  reg [63:0] out_data_R; // @[FPComputeNode.scala 66:27]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[FPComputeNode.scala 79:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[FPComputeNode.scala 85:27]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & left_valid_R; // @[FPComputeNode.scala 99:27]
  wire  _T_18 = _T_17 & right_valid_R; // @[FPComputeNode.scala 99:43]
  wire  _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire [14:0] _T_24 = value + 15'h1; // @[Counter.scala 39:22]
  wire  _T_26 = ~reset; // @[FPComputeNode.scala 108:17]
  wire [63:0] _T_19_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_16 = _T_18 ? _T_19_data : out_data_R; // @[FPComputeNode.scala 99:61]
  wire  _GEN_19 = _T_18 | out_valid_R_0; // @[FPComputeNode.scala 99:61]
  wire  _GEN_23 = _T_18 | state; // @[FPComputeNode.scala 99:61]
  wire  _T_29 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_45 = _T_16 & _T_18; // @[FPComputeNode.scala 108:17]
  FPUALU_1 FU ( // @[FPComputeNode.scala 64:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_16 ? _GEN_19 : out_valid_R_0; // @[HandShaking.scala 194:21 FPComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_16 : out_data_R; // @[FPComputeNode.scala 92:25 FPComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~left_valid_R; // @[FPComputeNode.scala 78:19]
  assign io_RightIO_ready = ~right_valid_R; // @[FPComputeNode.scala 84:20]
  assign FU_io_in1 = left_R_data; // @[FPComputeNode.scala 75:13]
  assign FU_io_in2 = right_R_data; // @[FPComputeNode.scala 76:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[14:0];
  _RAND_7 = {2{`RANDOM}};
  left_R_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  left_valid_R = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  right_R_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  task_ID_R = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_29) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_16) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_29) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        out_valid_R_0 <= _T_21;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      value <= 15'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        value <= _T_24;
      end
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= io_RightIO_bits_data;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_16) begin
      if (_T_18) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    task_ID_R <= enable_R_taskID;
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_23;
    end else if (state) begin
      if (_T_29) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_16) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_29) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_45 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [FPCompute] [FP_add2626] [Pred: %d] [Iter: %d] [In(0): %d] [In(1) %d] [Out: %d] [OpCode: fadd] [Cycle: %d]\n",task_ID_R,enable_R_control,value,left_R_data,right_R_data,FU_io_out,cycleCount); // @[FPComputeNode.scala 108:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStoreCache(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_SuccOp_0_ready,
  output        io_SuccOp_0_valid,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [63:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [63:0] io_inData_bits_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [63:0] io_MemReq_bits_addr,
  output [63:0] io_MemReq_bits_data,
  input         io_MemResp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 592:31]
  reg  enable_R_control; // @[HandShaking.scala 592:31]
  reg  enable_valid_R; // @[HandShaking.scala 593:31]
  reg  succ_ready_R_0; // @[HandShaking.scala 600:51]
  reg  succ_valid_R_0; // @[HandShaking.scala 601:51]
  wire  _T_5 = io_SuccOp_0_ready & io_SuccOp_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_5 ? 1'h0 : succ_valid_R_0; // @[HandShaking.scala 622:32]
  wire  _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_12 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [63:0] addr_R_data; // @[StoreCache.scala 59:23]
  reg [63:0] data_R_data; // @[StoreCache.scala 60:23]
  reg  addr_valid_R; // @[StoreCache.scala 61:29]
  reg  data_valid_R; // @[StoreCache.scala 62:29]
  reg [1:0] state; // @[StoreCache.scala 66:22]
  wire  _T_18 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_18 | addr_valid_R; // @[StoreCache.scala 80:27]
  wire  _T_19 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_19 | data_valid_R; // @[StoreCache.scala 85:26]
  wire  mem_req_fire = addr_valid_R & data_valid_R; // @[StoreCache.scala 102:51]
  wire  _T_38 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_40 = data_valid_R & addr_valid_R; // @[StoreCache.scala 154:27]
  wire  _T_41 = enable_R_control & mem_req_fire; // @[StoreCache.scala 155:33]
  wire  _GEN_28 = _T_40 & _T_41; // @[StoreCache.scala 154:44]
  wire  _GEN_33 = enable_valid_R & _GEN_28; // @[StoreCache.scala 153:51]
  wire  _T_44 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = io_MemResp_valid | _GEN_1; // @[StoreCache.scala 188:30]
  wire  _T_47 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_49 = &succ_ready_R_0; // @[HandShaking.scala 707:36]
  wire  _T_51 = &io_SuccOp_0_ready; // @[HandShaking.scala 707:72]
  wire  _T_52 = _T_49 | _T_51; // @[HandShaking.scala 707:41]
  wire [14:0] _T_62 = value + 15'h1; // @[Counter.scala 39:22]
  wire  _T_64 = ~reset; // @[StoreCache.scala 210:17]
  wire  _GEN_98 = ~_T_38; // @[StoreCache.scala 210:17]
  wire  _GEN_99 = ~_T_44; // @[StoreCache.scala 210:17]
  wire  _GEN_100 = _GEN_98 & _GEN_99; // @[StoreCache.scala 210:17]
  wire  _GEN_101 = _GEN_100 & _T_47; // @[StoreCache.scala 210:17]
  wire  _GEN_102 = _GEN_101 & _T_52; // @[StoreCache.scala 210:17]
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 650:19]
  assign io_SuccOp_0_valid = succ_valid_R_0; // @[HandShaking.scala 619:24]
  assign io_GepAddr_ready = ~addr_valid_R; // @[StoreCache.scala 75:20 StoreCache.scala 79:20]
  assign io_inData_ready = ~data_valid_R; // @[StoreCache.scala 76:19]
  assign io_MemReq_valid = _T_38 & _GEN_33; // @[StoreCache.scala 145:19 StoreCache.scala 156:29]
  assign io_MemReq_bits_addr = addr_R_data; // @[StoreCache.scala 139:23]
  assign io_MemReq_bits_data = data_R_data; // @[StoreCache.scala 140:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  succ_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  succ_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[14:0];
  _RAND_7 = {2{`RANDOM}};
  addr_R_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  data_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  data_valid_R = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_8) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_8) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_38) begin
      if (_T_8) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_44) begin
      if (_T_8) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_47) begin
      if (_T_52) begin
        enable_valid_R <= 1'h0;
      end else if (_T_8) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_8) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      succ_ready_R_0 <= 1'h0;
    end else if (_T_38) begin
      if (_T_5) begin
        succ_ready_R_0 <= io_SuccOp_0_ready;
      end
    end else if (_T_44) begin
      if (_T_5) begin
        succ_ready_R_0 <= io_SuccOp_0_ready;
      end
    end else if (_T_47) begin
      if (_T_52) begin
        succ_ready_R_0 <= 1'h0;
      end else if (_T_5) begin
        succ_ready_R_0 <= io_SuccOp_0_ready;
      end
    end else if (_T_5) begin
      succ_ready_R_0 <= io_SuccOp_0_ready;
    end
    if (reset) begin
      succ_valid_R_0 <= 1'h0;
    end else if (_T_38) begin
      if (enable_valid_R) begin
        if (_T_40) begin
          if (_T_41) begin
            if (_T_5) begin
              succ_valid_R_0 <= 1'h0;
            end
          end else begin
            succ_valid_R_0 <= 1'h1;
          end
        end else if (_T_5) begin
          succ_valid_R_0 <= 1'h0;
        end
      end else if (_T_5) begin
        succ_valid_R_0 <= 1'h0;
      end
    end else if (_T_44) begin
      succ_valid_R_0 <= _GEN_38;
    end else if (_T_5) begin
      succ_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_12;
    end
    if (reset) begin
      value <= 15'h0;
    end else if (!(_T_38)) begin
      if (!(_T_44)) begin
        if (_T_47) begin
          if (_T_52) begin
            value <= _T_62;
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_18) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_44) begin
      if (_T_18) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_47) begin
      if (_T_52) begin
        addr_R_data <= 64'h0;
      end else if (_T_18) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end else if (_T_18) begin
      addr_R_data <= io_GepAddr_bits_data;
    end
    if (reset) begin
      data_R_data <= 64'h0;
    end else if (_T_38) begin
      if (_T_19) begin
        data_R_data <= io_inData_bits_data;
      end
    end else if (_T_44) begin
      if (_T_19) begin
        data_R_data <= io_inData_bits_data;
      end
    end else if (_T_47) begin
      if (_T_52) begin
        data_R_data <= 64'h0;
      end else if (_T_19) begin
        data_R_data <= io_inData_bits_data;
      end
    end else if (_T_19) begin
      data_R_data <= io_inData_bits_data;
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else if (_T_38) begin
      addr_valid_R <= _GEN_13;
    end else if (_T_44) begin
      addr_valid_R <= _GEN_13;
    end else if (_T_47) begin
      if (_T_52) begin
        addr_valid_R <= 1'h0;
      end else begin
        addr_valid_R <= _GEN_13;
      end
    end else begin
      addr_valid_R <= _GEN_13;
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else if (_T_38) begin
      data_valid_R <= _GEN_17;
    end else if (_T_44) begin
      data_valid_R <= _GEN_17;
    end else if (_T_47) begin
      if (_T_52) begin
        data_valid_R <= 1'h0;
      end else begin
        data_valid_R <= _GEN_17;
      end
    end else begin
      data_valid_R <= _GEN_17;
    end
    if (reset) begin
      state <= 2'h0;
    end else if (_T_38) begin
      if (enable_valid_R) begin
        if (_T_40) begin
          if (_T_41) begin
            if (io_MemReq_ready) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end
    end else if (_T_44) begin
      if (io_MemResp_valid) begin
        state <= 2'h2;
      end
    end else if (_T_47) begin
      if (_T_52) begin
        state <= 2'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_102 & _T_64) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [STORE] [st_27] [Pred: %d] [Iter: %d] [Addr: %d] [Data: %d] [Cycle: %d]\n",enable_R_taskID,enable_R_control,value,addr_R_data,data_R_data,cycleCount); // @[StoreCache.scala 210:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_ready_R_1; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  reg  out_valid_R_1; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_8 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_13 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_15 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_23 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_29 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_30 = _T_29 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_36 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_37 = _T_2 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_39 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_32_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_19 = _T_30 ? _T_32_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_25 = _T_30 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_26 = _T_30 | out_valid_R_1; // @[ComputeNode.scala 147:81]
  wire  _GEN_31 = _T_30 | state; // @[ComputeNode.scala 147:81]
  wire  _T_43 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_44 = out_ready_R_1 | _T_2; // @[HandShaking.scala 251:83]
  wire  _T_45 = _T_43 & _T_44; // @[HandShaking.scala 252:27]
  wire  _GEN_62 = _T_23 & _T_30; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_23 ? _GEN_25 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_1_valid = _T_23 ? _GEN_26 : out_valid_R_1; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_1_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {2{`RANDOM}};
  left_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  right_R_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_4) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_4) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_45) begin
        enable_valid_R <= 1'h0;
      end else if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_4) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_2) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_0 <= _T_36;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_1 <= _T_37;
      end else if (_T_2) begin
        out_valid_R_1 <= 1'h0;
      end
    end else if (_T_2) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_8;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_13) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_13;
      end
    end else begin
      left_valid_R <= _GEN_13;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_15) begin
      right_R_data <= 64'h1;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_17;
      end
    end else begin
      right_valid_R <= _GEN_17;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_23) begin
      state <= _GEN_31;
    end else if (state) begin
      if (_T_45) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_23) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_45) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_indvars_iv_next28] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_10(
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out
);
  wire  _T_21 = io_in1 == io_in2; // @[Alu.scala 189:38]
  assign io_out = {{63'd0}, _T_21}; // @[Alu.scala 235:10]
endmodule
module ComputeNode_10(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_10 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h2;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [icmp_exitcond29] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: eq] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [63:0] io_CmpIO_bits_data,
  output        io_PredOp_0_ready,
  input         io_PredOp_0_valid,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1182:22]
  reg  cmp_R_control; // @[BranchNode.scala 1182:22]
  reg  cmp_valid; // @[BranchNode.scala 1183:26]
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1186:25]
  reg  enable_R_control; // @[BranchNode.scala 1186:25]
  reg  enable_valid_R; // @[BranchNode.scala 1187:31]
  reg  predecessor_valid_R_0; // @[BranchNode.scala 1191:61]
  reg  output_true_R_control; // @[BranchNode.scala 1193:30]
  reg  output_true_valid_R_0; // @[BranchNode.scala 1194:54]
  reg  fire_true_R_0; // @[BranchNode.scala 1195:46]
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1197:31]
  reg  output_false_R_control; // @[BranchNode.scala 1197:31]
  reg  output_false_valid_R_0; // @[BranchNode.scala 1198:56]
  reg  fire_false_R_0; // @[BranchNode.scala 1199:48]
  wire [4:0] task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1201:33]
  wire  _T_10 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = |io_CmpIO_bits_data; // @[BranchNode.scala 1207:44]
  wire  _GEN_4 = _T_10 | cmp_valid; // @[BranchNode.scala 1206:23]
  wire  _T_13 = io_PredOp_0_ready & io_PredOp_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_13 | predecessor_valid_R_0; // @[BranchNode.scala 1214:29]
  wire  _T_15 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = _T_15 | enable_valid_R; // @[BranchNode.scala 1232:24]
  wire  true_output = enable_R_control & cmp_R_control; // @[BranchNode.scala 1238:38]
  wire  _T_16 = ~cmp_R_control; // @[BranchNode.scala 1239:43]
  wire  false_output = enable_R_control & _T_16; // @[BranchNode.scala 1239:39]
  wire  _T_17 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_17 | fire_true_R_0; // @[BranchNode.scala 1250:33]
  wire  _GEN_14 = _T_17 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1250:33]
  wire  _T_18 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_18 | fire_false_R_0; // @[BranchNode.scala 1266:34]
  wire  _GEN_16 = _T_18 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1266:34]
  reg  state; // @[BranchNode.scala 1278:22]
  wire  _T_19 = ~state; // @[Conditional.scala 37:30]
  wire  _T_20 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1283:27]
  wire  _T_21 = _T_20 & predecessor_valid_R_0; // @[BranchNode.scala 1283:40]
  wire  _T_23 = ~reset; // @[BranchNode.scala 1293:21]
  wire  _GEN_17 = _T_21 | _GEN_14; // @[BranchNode.scala 1283:65]
  wire  _GEN_18 = _T_21 | _GEN_16; // @[BranchNode.scala 1283:65]
  wire  _GEN_19 = _T_21 | state; // @[BranchNode.scala 1283:65]
  wire  _T_29 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1313:27]
  wire  _GEN_80 = _T_19 & _T_21; // @[BranchNode.scala 1293:21]
  wire  _GEN_81 = _GEN_80 & enable_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_82 = _GEN_81 & cmp_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_86 = _GEN_81 & _T_16; // @[BranchNode.scala 1298:21]
  wire  _GEN_88 = ~enable_R_control; // @[BranchNode.scala 1304:19]
  wire  _GEN_89 = _GEN_80 & _GEN_88; // @[BranchNode.scala 1304:19]
  assign io_enable_ready = ~enable_valid_R; // @[BranchNode.scala 1231:19]
  assign io_CmpIO_ready = ~cmp_valid; // @[BranchNode.scala 1205:18]
  assign io_PredOp_0_ready = ~predecessor_valid_R_0; // @[BranchNode.scala 1213:24]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1246:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1245:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1262:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1261:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1261:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  predecessor_valid_R_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_true_R_control = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  output_false_R_control = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else if (_T_19) begin
      if (_T_10) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (state) begin
      if (_T_29) begin
        cmp_R_taskID <= 5'h0;
      end else if (_T_10) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (_T_10) begin
      cmp_R_taskID <= io_CmpIO_bits_taskID;
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else if (_T_19) begin
      if (_T_10) begin
        cmp_R_control <= _T_11;
      end
    end else if (state) begin
      if (_T_29) begin
        cmp_R_control <= 1'h0;
      end else if (_T_10) begin
        cmp_R_control <= _T_11;
      end
    end else if (_T_10) begin
      cmp_R_control <= _T_11;
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else if (_T_19) begin
      cmp_valid <= _GEN_4;
    end else if (state) begin
      if (_T_29) begin
        cmp_valid <= 1'h0;
      end else begin
        cmp_valid <= _GEN_4;
      end
    end else begin
      cmp_valid <= _GEN_4;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_19) begin
      if (_T_15) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_29) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_15) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_15) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_19) begin
      if (_T_15) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_29) begin
        enable_R_control <= 1'h0;
      end else if (_T_15) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_15) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_19) begin
      enable_valid_R <= _GEN_12;
    end else if (state) begin
      if (_T_29) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_12;
      end
    end else begin
      enable_valid_R <= _GEN_12;
    end
    if (reset) begin
      predecessor_valid_R_0 <= 1'h0;
    end else if (_T_19) begin
      predecessor_valid_R_0 <= _GEN_8;
    end else if (state) begin
      if (_T_29) begin
        predecessor_valid_R_0 <= 1'h0;
      end else begin
        predecessor_valid_R_0 <= _GEN_8;
      end
    end else begin
      predecessor_valid_R_0 <= _GEN_8;
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else if (_T_19) begin
      output_true_R_control <= true_output;
    end else if (state) begin
      if (_T_29) begin
        output_true_R_control <= 1'h0;
      end else begin
        output_true_R_control <= true_output;
      end
    end else begin
      output_true_R_control <= true_output;
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else if (_T_19) begin
      output_true_valid_R_0 <= _GEN_17;
    end else if (state) begin
      if (_T_29) begin
        output_true_valid_R_0 <= 1'h0;
      end else if (_T_17) begin
        output_true_valid_R_0 <= 1'h0;
      end
    end else if (_T_17) begin
      output_true_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else if (_T_19) begin
      fire_true_R_0 <= _GEN_13;
    end else if (state) begin
      if (_T_29) begin
        fire_true_R_0 <= 1'h0;
      end else begin
        fire_true_R_0 <= _GEN_13;
      end
    end else begin
      fire_true_R_0 <= _GEN_13;
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else if (_T_19) begin
      output_false_R_taskID <= task_id;
    end else if (state) begin
      if (_T_29) begin
        output_false_R_taskID <= 5'h0;
      end else begin
        output_false_R_taskID <= task_id;
      end
    end else begin
      output_false_R_taskID <= task_id;
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else if (_T_19) begin
      output_false_R_control <= false_output;
    end else if (state) begin
      if (_T_29) begin
        output_false_R_control <= 1'h0;
      end else begin
        output_false_R_control <= false_output;
      end
    end else begin
      output_false_R_control <= false_output;
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else if (_T_19) begin
      output_false_valid_R_0 <= _GEN_18;
    end else if (state) begin
      if (_T_29) begin
        output_false_valid_R_0 <= 1'h0;
      end else if (_T_18) begin
        output_false_valid_R_0 <= 1'h0;
      end
    end else if (_T_18) begin
      output_false_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else if (_T_19) begin
      fire_false_R_0 <= _GEN_15;
    end else if (state) begin
      if (_T_29) begin
        fire_false_R_0 <= 1'h0;
      end else begin
        fire_false_R_0 <= _GEN_15;
      end
    end else begin
      fire_false_R_0 <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_19) begin
      state <= _GEN_19;
    end else if (state) begin
      if (_T_29) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_30] [Out: T:1 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1293:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_86 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_30] [Out: T:0 - F:1] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1298:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_89 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_30] [Out: T:0 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1304:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_11(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_ready_R_1; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  reg  out_valid_R_1; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_8 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_13 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_15 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_23 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_29 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_30 = _T_29 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_36 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_37 = _T_2 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_39 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_32_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_19 = _T_30 ? _T_32_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_25 = _T_30 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_26 = _T_30 | out_valid_R_1; // @[ComputeNode.scala 147:81]
  wire  _GEN_31 = _T_30 | state; // @[ComputeNode.scala 147:81]
  wire  _T_43 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_44 = out_ready_R_1 | _T_2; // @[HandShaking.scala 251:83]
  wire  _T_45 = _T_43 & _T_44; // @[HandShaking.scala 252:27]
  wire  _GEN_62 = _T_23 & _T_30; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_23 ? _GEN_25 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_1_valid = _T_23 ? _GEN_26 : out_valid_R_1; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_1_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {2{`RANDOM}};
  left_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  right_R_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_4) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_4) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_45) begin
        enable_valid_R <= 1'h0;
      end else if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_4) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_2) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_0 <= _T_36;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_1 <= _T_37;
      end else if (_T_2) begin
        out_valid_R_1 <= 1'h0;
      end
    end else if (_T_2) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_8;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_13) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_13;
      end
    end else begin
      left_valid_R <= _GEN_13;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_15) begin
      right_R_data <= 64'h1;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_17;
      end
    end else begin
      right_valid_R <= _GEN_17;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_23) begin
      state <= _GEN_31;
    end else if (state) begin
      if (_T_45) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_23) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_45) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_indvars_iv_next7231] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_12(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_10 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h2;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [icmp_exitcond7732] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: eq] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [63:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1182:22]
  reg  cmp_R_control; // @[BranchNode.scala 1182:22]
  reg  cmp_valid; // @[BranchNode.scala 1183:26]
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1186:25]
  reg  enable_R_control; // @[BranchNode.scala 1186:25]
  reg  enable_valid_R; // @[BranchNode.scala 1187:31]
  reg  output_true_R_control; // @[BranchNode.scala 1193:30]
  reg  output_true_valid_R_0; // @[BranchNode.scala 1194:54]
  reg  fire_true_R_0; // @[BranchNode.scala 1195:46]
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1197:31]
  reg  output_false_R_control; // @[BranchNode.scala 1197:31]
  reg  output_false_valid_R_0; // @[BranchNode.scala 1198:56]
  reg  fire_false_R_0; // @[BranchNode.scala 1199:48]
  wire [4:0] task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1201:33]
  wire  _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  wire  _T_10 = |io_CmpIO_bits_data; // @[BranchNode.scala 1207:44]
  wire  _GEN_4 = _T_9 | cmp_valid; // @[BranchNode.scala 1206:23]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_12 | enable_valid_R; // @[BranchNode.scala 1232:24]
  wire  true_output = enable_R_control & cmp_R_control; // @[BranchNode.scala 1238:38]
  wire  _T_13 = ~cmp_R_control; // @[BranchNode.scala 1239:43]
  wire  false_output = enable_R_control & _T_13; // @[BranchNode.scala 1239:39]
  wire  _T_14 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_14 | fire_true_R_0; // @[BranchNode.scala 1250:33]
  wire  _GEN_10 = _T_14 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1250:33]
  wire  _T_15 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_15 | fire_false_R_0; // @[BranchNode.scala 1266:34]
  wire  _GEN_12 = _T_15 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1266:34]
  reg  state; // @[BranchNode.scala 1278:22]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1283:27]
  wire  _T_20 = ~reset; // @[BranchNode.scala 1293:21]
  wire  _GEN_13 = _T_17 | _GEN_10; // @[BranchNode.scala 1283:65]
  wire  _GEN_14 = _T_17 | _GEN_12; // @[BranchNode.scala 1283:65]
  wire  _GEN_15 = _T_17 | state; // @[BranchNode.scala 1283:65]
  wire  _T_26 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1313:27]
  wire  _GEN_73 = _T_16 & _T_17; // @[BranchNode.scala 1293:21]
  wire  _GEN_74 = _GEN_73 & enable_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_75 = _GEN_74 & cmp_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_79 = _GEN_74 & _T_13; // @[BranchNode.scala 1298:21]
  wire  _GEN_81 = ~enable_R_control; // @[BranchNode.scala 1304:19]
  wire  _GEN_82 = _GEN_73 & _GEN_81; // @[BranchNode.scala 1304:19]
  assign io_enable_ready = ~enable_valid_R; // @[BranchNode.scala 1231:19]
  assign io_CmpIO_ready = ~cmp_valid; // @[BranchNode.scala 1205:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1246:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1245:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1262:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1261:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1261:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_taskID <= 5'h0;
      end else if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (_T_9) begin
      cmp_R_taskID <= io_CmpIO_bits_taskID;
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_control <= 1'h0;
      end else if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (_T_9) begin
      cmp_R_control <= _T_10;
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else if (_T_16) begin
      cmp_valid <= _GEN_4;
    end else if (state) begin
      if (_T_26) begin
        cmp_valid <= 1'h0;
      end else begin
        cmp_valid <= _GEN_4;
      end
    end else begin
      cmp_valid <= _GEN_4;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_12) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      enable_valid_R <= _GEN_8;
    end else if (state) begin
      if (_T_26) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_8;
      end
    end else begin
      enable_valid_R <= _GEN_8;
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else if (_T_16) begin
      output_true_R_control <= true_output;
    end else if (state) begin
      if (_T_26) begin
        output_true_R_control <= 1'h0;
      end else begin
        output_true_R_control <= true_output;
      end
    end else begin
      output_true_R_control <= true_output;
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_true_valid_R_0 <= _GEN_13;
    end else if (state) begin
      if (_T_26) begin
        output_true_valid_R_0 <= 1'h0;
      end else if (_T_14) begin
        output_true_valid_R_0 <= 1'h0;
      end
    end else if (_T_14) begin
      output_true_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_true_R_0 <= _GEN_9;
    end else if (state) begin
      if (_T_26) begin
        fire_true_R_0 <= 1'h0;
      end else begin
        fire_true_R_0 <= _GEN_9;
      end
    end else begin
      fire_true_R_0 <= _GEN_9;
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else if (_T_16) begin
      output_false_R_taskID <= task_id;
    end else if (state) begin
      if (_T_26) begin
        output_false_R_taskID <= 5'h0;
      end else begin
        output_false_R_taskID <= task_id;
      end
    end else begin
      output_false_R_taskID <= task_id;
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else if (_T_16) begin
      output_false_R_control <= false_output;
    end else if (state) begin
      if (_T_26) begin
        output_false_R_control <= 1'h0;
      end else begin
        output_false_R_control <= false_output;
      end
    end else begin
      output_false_R_control <= false_output;
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_false_valid_R_0 <= _GEN_14;
    end else if (state) begin
      if (_T_26) begin
        output_false_valid_R_0 <= 1'h0;
      end else if (_T_15) begin
        output_false_valid_R_0 <= 1'h0;
      end
    end else if (_T_15) begin
      output_false_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_false_R_0 <= _GEN_11;
    end else if (state) begin
      if (_T_26) begin
        fire_false_R_0 <= 1'h0;
      end else begin
        fire_false_R_0 <= _GEN_11;
      end
    end else begin
      fire_false_R_0 <= _GEN_11;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_15;
    end else if (state) begin
      if (_T_26) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_33] [Out: T:1 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1293:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_33] [Out: T:0 - F:1] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1298:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_33] [Out: T:0 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1304:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_13(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_ready_R_1; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  reg  out_valid_R_1; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_8 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_13 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_15 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_23 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_29 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_30 = _T_29 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_36 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_37 = _T_2 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_39 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_32_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_19 = _T_30 ? _T_32_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_25 = _T_30 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_26 = _T_30 | out_valid_R_1; // @[ComputeNode.scala 147:81]
  wire  _GEN_31 = _T_30 | state; // @[ComputeNode.scala 147:81]
  wire  _T_43 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_44 = out_ready_R_1 | _T_2; // @[HandShaking.scala 251:83]
  wire  _T_45 = _T_43 & _T_44; // @[HandShaking.scala 252:27]
  wire  _GEN_62 = _T_23 & _T_30; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_23 ? _GEN_25 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_1_valid = _T_23 ? _GEN_26 : out_valid_R_1; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_1_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {2{`RANDOM}};
  left_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  right_R_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_4) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_4) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_45) begin
        enable_valid_R <= 1'h0;
      end else if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_4) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_2) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_0 <= _T_36;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_1 <= _T_37;
      end else if (_T_2) begin
        out_valid_R_1 <= 1'h0;
      end
    end else if (_T_2) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_8;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_13) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_13;
      end
    end else begin
      left_valid_R <= _GEN_13;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_15) begin
      right_R_data <= 64'h1;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_17;
      end
    end else begin
      right_valid_R <= _GEN_17;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_23) begin
      state <= _GEN_31;
    end else if (state) begin
      if (_T_45) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_23) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_45) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_indvars_iv_next7934] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_14(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_10 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h10;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [icmp_exitcond8135] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: eq] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [63:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1182:22]
  reg  cmp_R_control; // @[BranchNode.scala 1182:22]
  reg  cmp_valid; // @[BranchNode.scala 1183:26]
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1186:25]
  reg  enable_R_control; // @[BranchNode.scala 1186:25]
  reg  enable_valid_R; // @[BranchNode.scala 1187:31]
  reg  output_true_R_control; // @[BranchNode.scala 1193:30]
  reg  output_true_valid_R_0; // @[BranchNode.scala 1194:54]
  reg  fire_true_R_0; // @[BranchNode.scala 1195:46]
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1197:31]
  reg  output_false_R_control; // @[BranchNode.scala 1197:31]
  reg  output_false_valid_R_0; // @[BranchNode.scala 1198:56]
  reg  fire_false_R_0; // @[BranchNode.scala 1199:48]
  wire [4:0] task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1201:33]
  wire  _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  wire  _T_10 = |io_CmpIO_bits_data; // @[BranchNode.scala 1207:44]
  wire  _GEN_4 = _T_9 | cmp_valid; // @[BranchNode.scala 1206:23]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_12 | enable_valid_R; // @[BranchNode.scala 1232:24]
  wire  true_output = enable_R_control & cmp_R_control; // @[BranchNode.scala 1238:38]
  wire  _T_13 = ~cmp_R_control; // @[BranchNode.scala 1239:43]
  wire  false_output = enable_R_control & _T_13; // @[BranchNode.scala 1239:39]
  wire  _T_14 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_14 | fire_true_R_0; // @[BranchNode.scala 1250:33]
  wire  _GEN_10 = _T_14 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1250:33]
  wire  _T_15 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_15 | fire_false_R_0; // @[BranchNode.scala 1266:34]
  wire  _GEN_12 = _T_15 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1266:34]
  reg  state; // @[BranchNode.scala 1278:22]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1283:27]
  wire  _T_20 = ~reset; // @[BranchNode.scala 1293:21]
  wire  _GEN_13 = _T_17 | _GEN_10; // @[BranchNode.scala 1283:65]
  wire  _GEN_14 = _T_17 | _GEN_12; // @[BranchNode.scala 1283:65]
  wire  _GEN_15 = _T_17 | state; // @[BranchNode.scala 1283:65]
  wire  _T_26 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1313:27]
  wire  _GEN_73 = _T_16 & _T_17; // @[BranchNode.scala 1293:21]
  wire  _GEN_74 = _GEN_73 & enable_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_75 = _GEN_74 & cmp_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_79 = _GEN_74 & _T_13; // @[BranchNode.scala 1298:21]
  wire  _GEN_81 = ~enable_R_control; // @[BranchNode.scala 1304:19]
  wire  _GEN_82 = _GEN_73 & _GEN_81; // @[BranchNode.scala 1304:19]
  assign io_enable_ready = ~enable_valid_R; // @[BranchNode.scala 1231:19]
  assign io_CmpIO_ready = ~cmp_valid; // @[BranchNode.scala 1205:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1246:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1245:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1262:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1261:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1261:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_taskID <= 5'h0;
      end else if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (_T_9) begin
      cmp_R_taskID <= io_CmpIO_bits_taskID;
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_control <= 1'h0;
      end else if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (_T_9) begin
      cmp_R_control <= _T_10;
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else if (_T_16) begin
      cmp_valid <= _GEN_4;
    end else if (state) begin
      if (_T_26) begin
        cmp_valid <= 1'h0;
      end else begin
        cmp_valid <= _GEN_4;
      end
    end else begin
      cmp_valid <= _GEN_4;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_12) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      enable_valid_R <= _GEN_8;
    end else if (state) begin
      if (_T_26) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_8;
      end
    end else begin
      enable_valid_R <= _GEN_8;
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else if (_T_16) begin
      output_true_R_control <= true_output;
    end else if (state) begin
      if (_T_26) begin
        output_true_R_control <= 1'h0;
      end else begin
        output_true_R_control <= true_output;
      end
    end else begin
      output_true_R_control <= true_output;
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_true_valid_R_0 <= _GEN_13;
    end else if (state) begin
      if (_T_26) begin
        output_true_valid_R_0 <= 1'h0;
      end else if (_T_14) begin
        output_true_valid_R_0 <= 1'h0;
      end
    end else if (_T_14) begin
      output_true_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_true_R_0 <= _GEN_9;
    end else if (state) begin
      if (_T_26) begin
        fire_true_R_0 <= 1'h0;
      end else begin
        fire_true_R_0 <= _GEN_9;
      end
    end else begin
      fire_true_R_0 <= _GEN_9;
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else if (_T_16) begin
      output_false_R_taskID <= task_id;
    end else if (state) begin
      if (_T_26) begin
        output_false_R_taskID <= 5'h0;
      end else begin
        output_false_R_taskID <= task_id;
      end
    end else begin
      output_false_R_taskID <= task_id;
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else if (_T_16) begin
      output_false_R_control <= false_output;
    end else if (state) begin
      if (_T_26) begin
        output_false_R_control <= 1'h0;
      end else begin
        output_false_R_control <= false_output;
      end
    end else begin
      output_false_R_control <= false_output;
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_false_valid_R_0 <= _GEN_14;
    end else if (state) begin
      if (_T_26) begin
        output_false_valid_R_0 <= 1'h0;
      end else if (_T_15) begin
        output_false_valid_R_0 <= 1'h0;
      end
    end else if (_T_15) begin
      output_false_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_false_R_0 <= _GEN_11;
    end else if (state) begin
      if (_T_26) begin
        fire_false_R_0 <= 1'h0;
      end else begin
        fire_false_R_0 <= _GEN_11;
      end
    end else begin
      fire_false_R_0 <= _GEN_11;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_15;
    end else if (state) begin
      if (_T_26) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_36] [Out: T:1 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1293:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_36] [Out: T:0 - F:1] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1298:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_36] [Out: T:0 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1304:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_15(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_ready_R_1; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  reg  out_valid_R_1; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_8 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_13 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_15 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_23 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_29 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_30 = _T_29 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_36 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_37 = _T_2 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_39 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_32_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_19 = _T_30 ? _T_32_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_25 = _T_30 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_26 = _T_30 | out_valid_R_1; // @[ComputeNode.scala 147:81]
  wire  _GEN_31 = _T_30 | state; // @[ComputeNode.scala 147:81]
  wire  _T_43 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_44 = out_ready_R_1 | _T_2; // @[HandShaking.scala 251:83]
  wire  _T_45 = _T_43 & _T_44; // @[HandShaking.scala 252:27]
  wire  _GEN_62 = _T_23 & _T_30; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_23 ? _GEN_25 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_1_valid = _T_23 ? _GEN_26 : out_valid_R_1; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_1_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {2{`RANDOM}};
  left_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  right_R_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_4) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_4) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_45) begin
        enable_valid_R <= 1'h0;
      end else if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_4) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_2) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_0 <= _T_36;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_1 <= _T_37;
      end else if (_T_2) begin
        out_valid_R_1 <= 1'h0;
      end
    end else if (_T_2) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_8;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_13) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_13;
      end
    end else begin
      left_valid_R <= _GEN_13;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_15) begin
      right_R_data <= 64'h2;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_17;
      end
    end else begin
      right_valid_R <= _GEN_17;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_23) begin
      state <= _GEN_31;
    end else if (state) begin
      if (_T_45) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_23) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_45) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_indvars_iv_next8337] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_16(
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_out
);
  wire  _T_19 = io_in1 < io_in2; // @[Alu.scala 187:38]
  assign io_out = {{63'd0}, _T_19}; // @[Alu.scala 235:10]
endmodule
module ComputeNode_16(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_16 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h10;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [icmp_cmp238] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: slt] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [63:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output [4:0]  io_TrueOutput_0_bits_taskID,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output        io_FalseOutput_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1182:22]
  reg  cmp_R_control; // @[BranchNode.scala 1182:22]
  reg  cmp_valid; // @[BranchNode.scala 1183:26]
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1186:25]
  reg  enable_R_control; // @[BranchNode.scala 1186:25]
  reg  enable_valid_R; // @[BranchNode.scala 1187:31]
  reg [4:0] output_true_R_taskID; // @[BranchNode.scala 1193:30]
  reg  output_true_R_control; // @[BranchNode.scala 1193:30]
  reg  output_true_valid_R_0; // @[BranchNode.scala 1194:54]
  reg  fire_true_R_0; // @[BranchNode.scala 1195:46]
  reg  output_false_R_control; // @[BranchNode.scala 1197:31]
  reg  output_false_valid_R_0; // @[BranchNode.scala 1198:56]
  reg  fire_false_R_0; // @[BranchNode.scala 1199:48]
  wire [4:0] task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1201:33]
  wire  _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  wire  _T_10 = |io_CmpIO_bits_data; // @[BranchNode.scala 1207:44]
  wire  _GEN_4 = _T_9 | cmp_valid; // @[BranchNode.scala 1206:23]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_12 | enable_valid_R; // @[BranchNode.scala 1232:24]
  wire  true_output = enable_R_control & cmp_R_control; // @[BranchNode.scala 1238:38]
  wire  _T_13 = ~cmp_R_control; // @[BranchNode.scala 1239:43]
  wire  false_output = enable_R_control & _T_13; // @[BranchNode.scala 1239:39]
  wire  _T_14 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_14 | fire_true_R_0; // @[BranchNode.scala 1250:33]
  wire  _GEN_10 = _T_14 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1250:33]
  wire  _T_15 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_15 | fire_false_R_0; // @[BranchNode.scala 1266:34]
  wire  _GEN_12 = _T_15 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1266:34]
  reg  state; // @[BranchNode.scala 1278:22]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1283:27]
  wire  _T_20 = ~reset; // @[BranchNode.scala 1293:21]
  wire  _GEN_13 = _T_17 | _GEN_10; // @[BranchNode.scala 1283:65]
  wire  _GEN_14 = _T_17 | _GEN_12; // @[BranchNode.scala 1283:65]
  wire  _GEN_15 = _T_17 | state; // @[BranchNode.scala 1283:65]
  wire  _T_26 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1313:27]
  wire  _GEN_73 = _T_16 & _T_17; // @[BranchNode.scala 1293:21]
  wire  _GEN_74 = _GEN_73 & enable_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_75 = _GEN_74 & cmp_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_79 = _GEN_74 & _T_13; // @[BranchNode.scala 1298:21]
  wire  _GEN_81 = ~enable_R_control; // @[BranchNode.scala 1304:19]
  wire  _GEN_82 = _GEN_73 & _GEN_81; // @[BranchNode.scala 1304:19]
  assign io_enable_ready = ~enable_valid_R; // @[BranchNode.scala 1231:19]
  assign io_CmpIO_ready = ~cmp_valid; // @[BranchNode.scala 1205:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1246:28]
  assign io_TrueOutput_0_bits_taskID = output_true_R_taskID; // @[BranchNode.scala 1245:27]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1245:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1262:29]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1261:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_true_R_taskID = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  output_true_R_control = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_taskID <= 5'h0;
      end else if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (_T_9) begin
      cmp_R_taskID <= io_CmpIO_bits_taskID;
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_control <= 1'h0;
      end else if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (_T_9) begin
      cmp_R_control <= _T_10;
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else if (_T_16) begin
      cmp_valid <= _GEN_4;
    end else if (state) begin
      if (_T_26) begin
        cmp_valid <= 1'h0;
      end else begin
        cmp_valid <= _GEN_4;
      end
    end else begin
      cmp_valid <= _GEN_4;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_12) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      enable_valid_R <= _GEN_8;
    end else if (state) begin
      if (_T_26) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_8;
      end
    end else begin
      enable_valid_R <= _GEN_8;
    end
    if (reset) begin
      output_true_R_taskID <= 5'h0;
    end else if (_T_16) begin
      output_true_R_taskID <= task_id;
    end else if (state) begin
      if (_T_26) begin
        output_true_R_taskID <= 5'h0;
      end else begin
        output_true_R_taskID <= task_id;
      end
    end else begin
      output_true_R_taskID <= task_id;
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else if (_T_16) begin
      output_true_R_control <= true_output;
    end else if (state) begin
      if (_T_26) begin
        output_true_R_control <= 1'h0;
      end else begin
        output_true_R_control <= true_output;
      end
    end else begin
      output_true_R_control <= true_output;
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_true_valid_R_0 <= _GEN_13;
    end else if (state) begin
      if (_T_26) begin
        output_true_valid_R_0 <= 1'h0;
      end else if (_T_14) begin
        output_true_valid_R_0 <= 1'h0;
      end
    end else if (_T_14) begin
      output_true_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_true_R_0 <= _GEN_9;
    end else if (state) begin
      if (_T_26) begin
        fire_true_R_0 <= 1'h0;
      end else begin
        fire_true_R_0 <= _GEN_9;
      end
    end else begin
      fire_true_R_0 <= _GEN_9;
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else if (_T_16) begin
      output_false_R_control <= false_output;
    end else if (state) begin
      if (_T_26) begin
        output_false_R_control <= 1'h0;
      end else begin
        output_false_R_control <= false_output;
      end
    end else begin
      output_false_R_control <= false_output;
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_false_valid_R_0 <= _GEN_14;
    end else if (state) begin
      if (_T_26) begin
        output_false_valid_R_0 <= 1'h0;
      end else if (_T_15) begin
        output_false_valid_R_0 <= 1'h0;
      end
    end else if (_T_15) begin
      output_false_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_false_R_0 <= _GEN_11;
    end else if (state) begin
      if (_T_26) begin
        fire_false_R_0 <= 1'h0;
      end else begin
        fire_false_R_0 <= _GEN_11;
      end
    end else begin
      fire_false_R_0 <= _GEN_11;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_15;
    end else if (state) begin
      if (_T_26) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_39] [Out: T:1 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1293:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_39] [Out: T:0 - F:1] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1298:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_39] [Out: T:0 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1304:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_17(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [63:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_ready_R_1; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  reg  out_valid_R_1; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  wire  _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_8 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_13 = _T_13 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_17 = _T_15 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_23 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_29 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_30 = _T_29 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_36 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_37 = _T_2 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_39 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_32_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_19 = _T_30 ? _T_32_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_25 = _T_30 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_26 = _T_30 | out_valid_R_1; // @[ComputeNode.scala 147:81]
  wire  _GEN_31 = _T_30 | state; // @[ComputeNode.scala 147:81]
  wire  _T_43 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _T_44 = out_ready_R_1 | _T_2; // @[HandShaking.scala 251:83]
  wire  _T_45 = _T_43 & _T_44; // @[HandShaking.scala 252:27]
  wire  _GEN_62 = _T_23 & _T_30; // @[ComputeNode.scala 178:17]
  UALU_1 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_23 ? _GEN_25 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_1_valid = _T_23 ? _GEN_26 : out_valid_R_1; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_1_bits_data = _T_23 ? _GEN_19 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cycleCount = _RAND_7[14:0];
  _RAND_8 = {2{`RANDOM}};
  left_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  right_R_data = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  out_data_R = _RAND_13[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_4) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_4) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_45) begin
        enable_valid_R <= 1'h0;
      end else if (_T_4) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_4) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (state) begin
      if (_T_45) begin
        out_ready_R_1 <= 1'h0;
      end else if (_T_2) begin
        out_ready_R_1 <= io_Out_1_ready;
      end
    end else if (_T_2) begin
      out_ready_R_1 <= io_Out_1_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_0 <= _T_36;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        out_valid_R_1 <= _T_37;
      end else if (_T_2) begin
        out_valid_R_1 <= 1'h0;
      end
    end else if (_T_2) begin
      out_valid_R_1 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_8;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_13) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_13;
      end
    end else begin
      left_valid_R <= _GEN_13;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_15) begin
      right_R_data <= 64'h2;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_23) begin
      if (_T_30) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_17;
      end
    end else begin
      right_valid_R <= _GEN_17;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_23) begin
      state <= _GEN_31;
    end else if (state) begin
      if (_T_45) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_23) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_45) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [binaryOp_indvars_iv_next8540] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: add] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_18(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [63:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [63:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] FU_io_in1; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_in2; // @[ComputeNode.scala 61:18]
  wire [63:0] FU_io_out; // @[ComputeNode.scala 61:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 181:31]
  reg  enable_R_control; // @[HandShaking.scala 181:31]
  reg  enable_valid_R; // @[HandShaking.scala 182:31]
  reg  out_ready_R_0; // @[HandShaking.scala 185:46]
  reg  out_valid_R_0; // @[HandShaking.scala 186:46]
  wire  _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_7 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [63:0] left_R_data; // @[ComputeNode.scala 53:23]
  reg  left_valid_R; // @[ComputeNode.scala 54:29]
  reg [63:0] right_R_data; // @[ComputeNode.scala 57:24]
  reg  right_valid_R; // @[ComputeNode.scala 58:30]
  reg  state; // @[ComputeNode.scala 64:22]
  reg [63:0] out_data_R; // @[ComputeNode.scala 89:27]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 91:19]
  wire  _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_12 | left_valid_R; // @[ComputeNode.scala 105:26]
  wire  _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_15 = _T_14 | right_valid_R; // @[ComputeNode.scala 111:27]
  wire  _T_22 = ~state; // @[ComputeNode.scala 75:67]
  wire  _T_27 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 147:27]
  wire  _T_28 = _T_27 & right_valid_R; // @[ComputeNode.scala 147:43]
  wire  _T_32 = _T_1 ^ 1'h1; // @[HandShaking.scala 274:72]
  wire  _T_34 = ~reset; // @[ComputeNode.scala 178:17]
  wire [63:0] _T_30_data = FU_io_out; // @[interfaces.scala 289:20 interfaces.scala 290:15]
  wire [63:0] _GEN_17 = _T_28 ? _T_30_data : out_data_R; // @[ComputeNode.scala 147:81]
  wire  _GEN_20 = _T_28 | out_valid_R_0; // @[ComputeNode.scala 147:81]
  wire  _GEN_24 = _T_28 | state; // @[ComputeNode.scala 147:81]
  wire  _T_37 = out_ready_R_0 | _T_1; // @[HandShaking.scala 251:83]
  wire  _GEN_47 = _T_22 & _T_28; // @[ComputeNode.scala 178:17]
  UALU_16 FU ( // @[ComputeNode.scala 61:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign io_enable_ready = ~enable_valid_R; // @[HandShaking.scala 205:19]
  assign io_Out_0_valid = _T_22 ? _GEN_20 : out_valid_R_0; // @[HandShaking.scala 194:21 ComputeNode.scala 172:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_Out_0_bits_data = _T_22 ? _GEN_17 : out_data_R; // @[ComputeNode.scala 137:25 ComputeNode.scala 170:33]
  assign io_LeftIO_ready = ~left_valid_R; // @[ComputeNode.scala 104:19]
  assign io_RightIO_ready = ~right_valid_R; // @[ComputeNode.scala 110:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 101:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 102:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cycleCount = _RAND_5[14:0];
  _RAND_6 = {2{`RANDOM}};
  left_R_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  right_R_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  out_data_R = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_3) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_3) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (state) begin
      if (_T_37) begin
        enable_valid_R <= 1'h0;
      end else if (_T_3) begin
        enable_valid_R <= io_enable_valid;
      end
    end else if (_T_3) begin
      enable_valid_R <= io_enable_valid;
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (state) begin
      if (_T_37) begin
        out_ready_R_0 <= 1'h0;
      end else if (_T_1) begin
        out_ready_R_0 <= io_Out_0_ready;
      end
    end else if (_T_1) begin
      out_ready_R_0 <= io_Out_0_ready;
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        out_valid_R_0 <= _T_32;
      end else if (_T_1) begin
        out_valid_R_0 <= 1'h0;
      end
    end else if (_T_1) begin
      out_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_7;
    end
    if (reset) begin
      left_R_data <= 64'h0;
    end else if (_T_12) begin
      left_R_data <= io_LeftIO_bits_data;
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        left_valid_R <= 1'h0;
      end else begin
        left_valid_R <= _GEN_11;
      end
    end else begin
      left_valid_R <= _GEN_11;
    end
    if (reset) begin
      right_R_data <= 64'h0;
    end else if (_T_14) begin
      right_R_data <= 64'h10;
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else if (_T_22) begin
      if (_T_28) begin
        right_valid_R <= 1'h0;
      end else begin
        right_valid_R <= _GEN_15;
      end
    end else begin
      right_valid_R <= _GEN_15;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_22) begin
      state <= _GEN_24;
    end else if (state) begin
      if (_T_37) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      out_data_R <= 64'h0;
    end else if (_T_22) begin
      if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (state) begin
      if (_T_37) begin
        out_data_R <= 64'h0;
      end else if (enable_R_control) begin
        out_data_R <= FU_io_out;
      end else begin
        out_data_R <= 64'h0;
      end
    end else if (enable_R_control) begin
      out_data_R <= FU_io_out;
    end else begin
      out_data_R <= 64'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_47 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [COMPUTE] [icmp_cmp41] [Pred: %d] [In(0): 0x%x] [In(1) 0x%x] [Out: 0x%x] [OpCode: slt] [Cycle: %d]\n",taskID,enable_R_control,left_R_data,right_R_data,FU_io_out,cycleCount); // @[ComputeNode.scala 178:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [63:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output [4:0]  io_TrueOutput_0_bits_taskID,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output        io_FalseOutput_0_bits_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1182:22]
  reg  cmp_R_control; // @[BranchNode.scala 1182:22]
  reg  cmp_valid; // @[BranchNode.scala 1183:26]
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1186:25]
  reg  enable_R_control; // @[BranchNode.scala 1186:25]
  reg  enable_valid_R; // @[BranchNode.scala 1187:31]
  reg [4:0] output_true_R_taskID; // @[BranchNode.scala 1193:30]
  reg  output_true_R_control; // @[BranchNode.scala 1193:30]
  reg  output_true_valid_R_0; // @[BranchNode.scala 1194:54]
  reg  fire_true_R_0; // @[BranchNode.scala 1195:46]
  reg  output_false_R_control; // @[BranchNode.scala 1197:31]
  reg  output_false_valid_R_0; // @[BranchNode.scala 1198:56]
  reg  fire_false_R_0; // @[BranchNode.scala 1199:48]
  wire [4:0] task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1201:33]
  wire  _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  wire  _T_10 = |io_CmpIO_bits_data; // @[BranchNode.scala 1207:44]
  wire  _GEN_4 = _T_9 | cmp_valid; // @[BranchNode.scala 1206:23]
  wire  _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_12 | enable_valid_R; // @[BranchNode.scala 1232:24]
  wire  true_output = enable_R_control & cmp_R_control; // @[BranchNode.scala 1238:38]
  wire  _T_13 = ~cmp_R_control; // @[BranchNode.scala 1239:43]
  wire  false_output = enable_R_control & _T_13; // @[BranchNode.scala 1239:39]
  wire  _T_14 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_9 = _T_14 | fire_true_R_0; // @[BranchNode.scala 1250:33]
  wire  _GEN_10 = _T_14 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1250:33]
  wire  _T_15 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_15 | fire_false_R_0; // @[BranchNode.scala 1266:34]
  wire  _GEN_12 = _T_15 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1266:34]
  reg  state; // @[BranchNode.scala 1278:22]
  wire  _T_16 = ~state; // @[Conditional.scala 37:30]
  wire  _T_17 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1283:27]
  wire  _T_20 = ~reset; // @[BranchNode.scala 1293:21]
  wire  _GEN_13 = _T_17 | _GEN_10; // @[BranchNode.scala 1283:65]
  wire  _GEN_14 = _T_17 | _GEN_12; // @[BranchNode.scala 1283:65]
  wire  _GEN_15 = _T_17 | state; // @[BranchNode.scala 1283:65]
  wire  _T_26 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1313:27]
  wire  _GEN_73 = _T_16 & _T_17; // @[BranchNode.scala 1293:21]
  wire  _GEN_74 = _GEN_73 & enable_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_75 = _GEN_74 & cmp_R_control; // @[BranchNode.scala 1293:21]
  wire  _GEN_79 = _GEN_74 & _T_13; // @[BranchNode.scala 1298:21]
  wire  _GEN_81 = ~enable_R_control; // @[BranchNode.scala 1304:19]
  wire  _GEN_82 = _GEN_73 & _GEN_81; // @[BranchNode.scala 1304:19]
  assign io_enable_ready = ~enable_valid_R; // @[BranchNode.scala 1231:19]
  assign io_CmpIO_ready = ~cmp_valid; // @[BranchNode.scala 1205:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1246:28]
  assign io_TrueOutput_0_bits_taskID = output_true_R_taskID; // @[BranchNode.scala 1245:27]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1245:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1262:29]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1261:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  output_true_R_taskID = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  output_true_R_control = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_taskID <= 5'h0;
      end else if (_T_9) begin
        cmp_R_taskID <= io_CmpIO_bits_taskID;
      end
    end else if (_T_9) begin
      cmp_R_taskID <= io_CmpIO_bits_taskID;
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (state) begin
      if (_T_26) begin
        cmp_R_control <= 1'h0;
      end else if (_T_9) begin
        cmp_R_control <= _T_10;
      end
    end else if (_T_9) begin
      cmp_R_control <= _T_10;
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else if (_T_16) begin
      cmp_valid <= _GEN_4;
    end else if (state) begin
      if (_T_26) begin
        cmp_valid <= 1'h0;
      end else begin
        cmp_valid <= _GEN_4;
      end
    end else begin
      cmp_valid <= _GEN_4;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_taskID <= 5'h0;
      end else if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end else if (_T_12) begin
      enable_R_taskID <= io_enable_bits_taskID;
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_16) begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (state) begin
      if (_T_26) begin
        enable_R_control <= 1'h0;
      end else if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end else if (_T_12) begin
      enable_R_control <= io_enable_bits_control;
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_16) begin
      enable_valid_R <= _GEN_8;
    end else if (state) begin
      if (_T_26) begin
        enable_valid_R <= 1'h0;
      end else begin
        enable_valid_R <= _GEN_8;
      end
    end else begin
      enable_valid_R <= _GEN_8;
    end
    if (reset) begin
      output_true_R_taskID <= 5'h0;
    end else if (_T_16) begin
      output_true_R_taskID <= task_id;
    end else if (state) begin
      if (_T_26) begin
        output_true_R_taskID <= 5'h0;
      end else begin
        output_true_R_taskID <= task_id;
      end
    end else begin
      output_true_R_taskID <= task_id;
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else if (_T_16) begin
      output_true_R_control <= true_output;
    end else if (state) begin
      if (_T_26) begin
        output_true_R_control <= 1'h0;
      end else begin
        output_true_R_control <= true_output;
      end
    end else begin
      output_true_R_control <= true_output;
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_true_valid_R_0 <= _GEN_13;
    end else if (state) begin
      if (_T_26) begin
        output_true_valid_R_0 <= 1'h0;
      end else if (_T_14) begin
        output_true_valid_R_0 <= 1'h0;
      end
    end else if (_T_14) begin
      output_true_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_true_R_0 <= _GEN_9;
    end else if (state) begin
      if (_T_26) begin
        fire_true_R_0 <= 1'h0;
      end else begin
        fire_true_R_0 <= _GEN_9;
      end
    end else begin
      fire_true_R_0 <= _GEN_9;
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else if (_T_16) begin
      output_false_R_control <= false_output;
    end else if (state) begin
      if (_T_26) begin
        output_false_R_control <= 1'h0;
      end else begin
        output_false_R_control <= false_output;
      end
    end else begin
      output_false_R_control <= false_output;
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else if (_T_16) begin
      output_false_valid_R_0 <= _GEN_14;
    end else if (state) begin
      if (_T_26) begin
        output_false_valid_R_0 <= 1'h0;
      end else if (_T_15) begin
        output_false_valid_R_0 <= 1'h0;
      end
    end else if (_T_15) begin
      output_false_valid_R_0 <= 1'h0;
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else if (_T_16) begin
      fire_false_R_0 <= _GEN_11;
    end else if (state) begin
      if (_T_26) begin
        fire_false_R_0 <= 1'h0;
      end else begin
        fire_false_R_0 <= _GEN_11;
      end
    end else begin
      fire_false_R_0 <= _GEN_11;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_16) begin
      state <= _GEN_15;
    end else if (state) begin
      if (_T_26) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_42] [Out: T:1 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1293:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_42] [Out: T:0 - F:1] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1298:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_82 & _T_20) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CBR] [br_42] [Out: T:0 - F:0] [Cycle: %d]\n",task_id,cycleCount); // @[BranchNode.scala 1304:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module RetNode2(
  input        clock,
  input        reset,
  output       io_In_enable_ready,
  input        io_In_enable_valid,
  input  [4:0] io_In_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg  state; // @[RetNode.scala 141:22]
  reg  enable_valid_R; // @[RetNode.scala 144:31]
  reg [4:0] output_R_enable_taskID; // @[RetNode.scala 150:25]
  reg  out_ready_R; // @[RetNode.scala 151:28]
  reg  out_valid_R; // @[RetNode.scala 152:28]
  wire  _T_6 = io_In_enable_ready & io_In_enable_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_7 ? 1'h0 : out_valid_R; // @[RetNode.scala 194:23]
  wire  _T_8 = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_11 = enable_valid_R | _GEN_8; // @[RetNode.scala 202:28]
  wire  _GEN_12 = enable_valid_R | state; // @[RetNode.scala 202:28]
  wire  _T_11 = ~reset; // @[RetNode.scala 221:17]
  wire  _GEN_25 = ~_T_8; // @[RetNode.scala 221:17]
  wire  _GEN_26 = _GEN_25 & state; // @[RetNode.scala 221:17]
  wire  _GEN_27 = _GEN_26 & out_ready_R; // @[RetNode.scala 221:17]
  assign io_In_enable_ready = ~enable_valid_R; // @[RetNode.scala 163:22]
  assign io_Out_valid = out_valid_R; // @[RetNode.scala 180:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  output_R_enable_taskID = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  out_ready_R = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  out_valid_R = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_8) begin
      state <= _GEN_12;
    end else if (state) begin
      if (out_ready_R) begin
        state <= 1'h0;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_8) begin
      if (_T_6) begin
        enable_valid_R <= io_In_enable_valid;
      end
    end else if (state) begin
      if (out_ready_R) begin
        enable_valid_R <= 1'h0;
      end else if (_T_6) begin
        enable_valid_R <= io_In_enable_valid;
      end
    end else if (_T_6) begin
      enable_valid_R <= io_In_enable_valid;
    end
    if (reset) begin
      output_R_enable_taskID <= 5'h0;
    end else if (_T_6) begin
      output_R_enable_taskID <= io_In_enable_bits_taskID;
    end
    if (reset) begin
      out_ready_R <= 1'h0;
    end else if (_T_8) begin
      if (_T_7) begin
        out_ready_R <= io_Out_ready;
      end
    end else if (state) begin
      if (out_ready_R) begin
        out_ready_R <= 1'h0;
      end else if (_T_7) begin
        out_ready_R <= io_Out_ready;
      end
    end else if (_T_7) begin
      out_ready_R <= io_Out_ready;
    end
    if (reset) begin
      out_valid_R <= 1'h0;
    end else if (_T_8) begin
      out_valid_R <= _GEN_11;
    end else if (state) begin
      if (out_ready_R) begin
        out_valid_R <= 1'h0;
      end else if (_T_7) begin
        out_valid_R <= 1'h0;
      end
    end else if (_T_7) begin
      out_valid_R <= 1'h0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_11) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [ret_43] [Cycle: %d]\n",output_R_enable_taskID,cycleCount); // @[RetNode.scala 221:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 113:25]
  reg  enable_R_control; // @[ConstNode.scala 113:25]
  reg  enable_valid_R; // @[ConstNode.scala 114:31]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 116:19]
  reg  state; // @[ConstNode.scala 135:22]
  wire  _T_7 = ~state; // @[Conditional.scala 37:30]
  wire  _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~reset; // @[ConstNode.scala 149:17]
  wire  _GEN_7 = _T_8 | enable_valid_R; // @[ConstNode.scala 139:30]
  wire  _GEN_29 = _T_7 & _T_8; // @[ConstNode.scala 149:17]
  assign io_enable_ready = ~enable_valid_R; // @[ConstNode.scala 126:19]
  assign io_Out_valid = _T_7 ? _GEN_7 : enable_valid_R; // @[ConstNode.scala 127:16 ConstNode.scala 140:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 129:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_taskID <= 5'h0;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_control <= io_enable_bits_control;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_control <= 1'h0;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_valid_R <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_valid_R <= 1'h0;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (_T_9) begin
          state <= 1'h0;
        end else begin
          state <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & _T_11) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CONST] [Bbgemm] [Pred: %d] [Val: 0x%x] [Cycle: %d]\n",taskID,enable_R_control,64'h0,cycleCount); // @[ConstNode.scala 149:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_3(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 113:25]
  reg  enable_R_control; // @[ConstNode.scala 113:25]
  reg  enable_valid_R; // @[ConstNode.scala 114:31]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 116:19]
  reg  state; // @[ConstNode.scala 135:22]
  wire  _T_7 = ~state; // @[Conditional.scala 37:30]
  wire  _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~reset; // @[ConstNode.scala 149:17]
  wire  _GEN_7 = _T_8 | enable_valid_R; // @[ConstNode.scala 139:30]
  wire  _GEN_29 = _T_7 & _T_8; // @[ConstNode.scala 149:17]
  assign io_enable_ready = ~enable_valid_R; // @[ConstNode.scala 126:19]
  assign io_Out_valid = _T_7 ? _GEN_7 : enable_valid_R; // @[ConstNode.scala 127:16 ConstNode.scala 140:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_taskID <= 5'h0;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_control <= io_enable_bits_control;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_control <= 1'h0;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_valid_R <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_valid_R <= 1'h0;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (_T_9) begin
          state <= 1'h0;
        end else begin
          state <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & _T_11) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CONST] [Bbgemm] [Pred: %d] [Val: 0x%x] [Cycle: %d]\n",taskID,enable_R_control,64'h4,cycleCount); // @[ConstNode.scala 149:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_7(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 113:25]
  reg  enable_R_control; // @[ConstNode.scala 113:25]
  reg  enable_valid_R; // @[ConstNode.scala 114:31]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 116:19]
  reg  state; // @[ConstNode.scala 135:22]
  wire  _T_7 = ~state; // @[Conditional.scala 37:30]
  wire  _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~reset; // @[ConstNode.scala 149:17]
  wire  _GEN_7 = _T_8 | enable_valid_R; // @[ConstNode.scala 139:30]
  wire  _GEN_29 = _T_7 & _T_8; // @[ConstNode.scala 149:17]
  assign io_enable_ready = ~enable_valid_R; // @[ConstNode.scala 126:19]
  assign io_Out_valid = _T_7 ? _GEN_7 : enable_valid_R; // @[ConstNode.scala 127:16 ConstNode.scala 140:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_taskID <= 5'h0;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_control <= io_enable_bits_control;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_control <= 1'h0;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_valid_R <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_valid_R <= 1'h0;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (_T_9) begin
          state <= 1'h0;
        end else begin
          state <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & _T_11) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CONST] [Bbgemm] [Pred: %d] [Val: 0x%x] [Cycle: %d]\n",taskID,enable_R_control,64'h1,cycleCount); // @[ConstNode.scala 149:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_8(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 113:25]
  reg  enable_R_control; // @[ConstNode.scala 113:25]
  reg  enable_valid_R; // @[ConstNode.scala 114:31]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 116:19]
  reg  state; // @[ConstNode.scala 135:22]
  wire  _T_7 = ~state; // @[Conditional.scala 37:30]
  wire  _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~reset; // @[ConstNode.scala 149:17]
  wire  _GEN_7 = _T_8 | enable_valid_R; // @[ConstNode.scala 139:30]
  wire  _GEN_29 = _T_7 & _T_8; // @[ConstNode.scala 149:17]
  assign io_enable_ready = ~enable_valid_R; // @[ConstNode.scala 126:19]
  assign io_Out_valid = _T_7 ? _GEN_7 : enable_valid_R; // @[ConstNode.scala 127:16 ConstNode.scala 140:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_taskID <= 5'h0;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_control <= io_enable_bits_control;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_control <= 1'h0;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_valid_R <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_valid_R <= 1'h0;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (_T_9) begin
          state <= 1'h0;
        end else begin
          state <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & _T_11) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CONST] [Bbgemm] [Pred: %d] [Val: 0x%x] [Cycle: %d]\n",taskID,enable_R_control,64'h2,cycleCount); // @[ConstNode.scala 149:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_12(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [14:0] cycleCount; // @[Counter.scala 29:33]
  wire [14:0] _T_3 = cycleCount + 15'h1; // @[Counter.scala 39:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 113:25]
  reg  enable_R_control; // @[ConstNode.scala 113:25]
  reg  enable_valid_R; // @[ConstNode.scala 114:31]
  wire [4:0] taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 116:19]
  reg  state; // @[ConstNode.scala 135:22]
  wire  _T_7 = ~state; // @[Conditional.scala 37:30]
  wire  _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  wire  _T_11 = ~reset; // @[ConstNode.scala 149:17]
  wire  _GEN_7 = _T_8 | enable_valid_R; // @[ConstNode.scala 139:30]
  wire  _GEN_29 = _T_7 & _T_8; // @[ConstNode.scala 149:17]
  assign io_enable_ready = ~enable_valid_R; // @[ConstNode.scala 126:19]
  assign io_Out_valid = _T_7 ? _GEN_7 : enable_valid_R; // @[ConstNode.scala 127:16 ConstNode.scala 140:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycleCount = _RAND_0[14:0];
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cycleCount <= 15'h0;
    end else begin
      cycleCount <= _T_3;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_taskID <= 5'h0;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_R_control <= io_enable_bits_control;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_R_control <= 1'h0;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (!(_T_9)) begin
          enable_valid_R <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        enable_valid_R <= 1'h0;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else if (_T_7) begin
      if (_T_8) begin
        if (_T_9) begin
          state <= 1'h0;
        end else begin
          state <= 1'h1;
        end
      end
    end else if (state) begin
      if (_T_9) begin
        state <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_29 & _T_11) begin
          $fwrite(32'h80000002,"[LOG] [Bbgemm] [TID: %d] [CONST] [Bbgemm] [Pred: %d] [Val: 0x%x] [Cycle: %d]\n",taskID,enable_R_control,64'h10,cycleCount); // @[ConstNode.scala 149:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module bbgemmDF(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_dataPtrs_field2_data,
  input  [31:0] io_in_bits_dataPtrs_field1_data,
  input  [31:0] io_in_bits_dataPtrs_field0_data,
  input         io_MemResp_valid,
  input  [63:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [63:0] io_MemReq_bits_addr,
  output [63:0] io_MemReq_bits_data,
  output [7:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  input         io_out_ready,
  output        io_out_valid
);
  wire  MemCtrl_clock; // @[bbgemm.scala 34:23]
  wire  MemCtrl_reset; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_0_MemReq_ready; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_0_MemReq_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_rd_mem_0_MemReq_bits_addr; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_0_MemResp_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_rd_mem_0_MemResp_bits_data; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_1_MemReq_ready; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_1_MemReq_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_rd_mem_1_MemReq_bits_addr; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_1_MemResp_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_rd_mem_1_MemResp_bits_data; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_2_MemReq_ready; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_2_MemReq_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_rd_mem_2_MemReq_bits_addr; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_rd_mem_2_MemResp_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_rd_mem_2_MemResp_bits_data; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_wr_mem_0_MemReq_ready; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_wr_mem_0_MemReq_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_wr_mem_0_MemReq_bits_addr; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_wr_mem_0_MemReq_bits_data; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_wr_mem_0_MemResp_valid; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_cache_MemReq_ready; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_cache_MemReq_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_cache_MemReq_bits_addr; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_cache_MemReq_bits_data; // @[bbgemm.scala 34:23]
  wire [7:0] MemCtrl_io_cache_MemReq_bits_mask; // @[bbgemm.scala 34:23]
  wire [7:0] MemCtrl_io_cache_MemReq_bits_tag; // @[bbgemm.scala 34:23]
  wire  MemCtrl_io_cache_MemResp_valid; // @[bbgemm.scala 34:23]
  wire [63:0] MemCtrl_io_cache_MemResp_bits_data; // @[bbgemm.scala 34:23]
  wire [7:0] MemCtrl_io_cache_MemResp_bits_tag; // @[bbgemm.scala 34:23]
  wire  ArgSplitter_clock; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_reset; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_In_ready; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_In_valid; // @[bbgemm.scala 38:27]
  wire [63:0] ArgSplitter_io_In_bits_dataPtrs_field2_data; // @[bbgemm.scala 38:27]
  wire [63:0] ArgSplitter_io_In_bits_dataPtrs_field1_data; // @[bbgemm.scala 38:27]
  wire [63:0] ArgSplitter_io_In_bits_dataPtrs_field0_data; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_enable_ready; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_enable_valid; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_enable_bits_control; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_dataPtrs_field2_0_ready; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_dataPtrs_field2_0_valid; // @[bbgemm.scala 38:27]
  wire [63:0] ArgSplitter_io_Out_dataPtrs_field2_0_bits_data; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_dataPtrs_field1_0_ready; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_dataPtrs_field1_0_valid; // @[bbgemm.scala 38:27]
  wire [63:0] ArgSplitter_io_Out_dataPtrs_field1_0_bits_data; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_dataPtrs_field0_0_ready; // @[bbgemm.scala 38:27]
  wire  ArgSplitter_io_Out_dataPtrs_field0_0_valid; // @[bbgemm.scala 38:27]
  wire [63:0] ArgSplitter_io_Out_dataPtrs_field0_0_bits_data; // @[bbgemm.scala 38:27]
  wire  Loop_0_clock; // @[bbgemm.scala 47:22]
  wire  Loop_0_reset; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_enable_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_enable_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_enable_bits_taskID; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_enable_bits_control; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_InLiveIn_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_1_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_1_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_InLiveIn_1_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_2_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_2_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_InLiveIn_2_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_3_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_3_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_InLiveIn_3_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_4_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_4_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_InLiveIn_4_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_5_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_InLiveIn_5_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_InLiveIn_5_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field5_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field5_1_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field5_1_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field5_1_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field4_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_activate_loop_start_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_activate_loop_start_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_activate_loop_start_bits_control; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_activate_loop_back_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_activate_loop_back_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_activate_loop_back_bits_control; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopBack_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopBack_0_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_loopBack_0_bits_taskID; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopBack_0_bits_control; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopFinish_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopFinish_0_valid; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopFinish_0_bits_control; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_CarryDepenIn_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_CarryDepenIn_0_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 47:22]
  wire [63:0] Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopExit_0_ready; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopExit_0_valid; // @[bbgemm.scala 47:22]
  wire [4:0] Loop_0_io_loopExit_0_bits_taskID; // @[bbgemm.scala 47:22]
  wire  Loop_0_io_loopExit_0_bits_control; // @[bbgemm.scala 47:22]
  wire  Loop_1_clock; // @[bbgemm.scala 49:22]
  wire  Loop_1_reset; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_enable_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_enable_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_enable_bits_taskID; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_enable_bits_control; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_InLiveIn_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_1_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_1_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_InLiveIn_1_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_2_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_2_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_InLiveIn_2_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_3_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_3_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_InLiveIn_3_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_4_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_4_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_InLiveIn_4_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_5_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_InLiveIn_5_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_InLiveIn_5_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field5_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field4_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field4_1_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field4_1_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field4_1_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field0_1_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_OutLiveIn_field0_1_valid; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_OutLiveIn_field0_1_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_activate_loop_start_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_activate_loop_start_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_activate_loop_start_bits_control; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_activate_loop_back_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_activate_loop_back_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_activate_loop_back_bits_control; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopBack_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopBack_0_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_loopBack_0_bits_taskID; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopBack_0_bits_control; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopFinish_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopFinish_0_valid; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopFinish_0_bits_control; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_CarryDepenIn_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_CarryDepenIn_0_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 49:22]
  wire [63:0] Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopExit_0_ready; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopExit_0_valid; // @[bbgemm.scala 49:22]
  wire [4:0] Loop_1_io_loopExit_0_bits_taskID; // @[bbgemm.scala 49:22]
  wire  Loop_1_io_loopExit_0_bits_control; // @[bbgemm.scala 49:22]
  wire  Loop_2_clock; // @[bbgemm.scala 51:22]
  wire  Loop_2_reset; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_enable_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_enable_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_enable_bits_taskID; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_enable_bits_control; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_0_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_InLiveIn_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_1_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_1_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_InLiveIn_1_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_2_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_2_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_InLiveIn_2_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_3_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_3_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_InLiveIn_3_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_4_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_InLiveIn_4_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_InLiveIn_4_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field4_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_activate_loop_start_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_activate_loop_start_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_activate_loop_start_bits_control; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_activate_loop_back_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_activate_loop_back_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_activate_loop_back_bits_control; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopBack_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopBack_0_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_loopBack_0_bits_taskID; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopBack_0_bits_control; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopFinish_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopFinish_0_valid; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopFinish_0_bits_control; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_CarryDepenIn_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_CarryDepenIn_0_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 51:22]
  wire [63:0] Loop_2_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopExit_0_ready; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopExit_0_valid; // @[bbgemm.scala 51:22]
  wire [4:0] Loop_2_io_loopExit_0_bits_taskID; // @[bbgemm.scala 51:22]
  wire  Loop_2_io_loopExit_0_bits_control; // @[bbgemm.scala 51:22]
  wire  Loop_3_clock; // @[bbgemm.scala 53:22]
  wire  Loop_3_reset; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_enable_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_enable_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_enable_bits_taskID; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_enable_bits_control; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_0_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_InLiveIn_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_1_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_1_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_InLiveIn_1_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_2_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_2_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_InLiveIn_2_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_3_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_InLiveIn_3_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_InLiveIn_3_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_activate_loop_start_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_activate_loop_start_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_activate_loop_start_bits_control; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_activate_loop_back_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_activate_loop_back_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_activate_loop_back_bits_control; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopBack_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopBack_0_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_loopBack_0_bits_taskID; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopBack_0_bits_control; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopFinish_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopFinish_0_valid; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopFinish_0_bits_control; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_CarryDepenIn_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_CarryDepenIn_0_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 53:22]
  wire [63:0] Loop_3_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopExit_0_ready; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopExit_0_valid; // @[bbgemm.scala 53:22]
  wire [4:0] Loop_3_io_loopExit_0_bits_taskID; // @[bbgemm.scala 53:22]
  wire  Loop_3_io_loopExit_0_bits_control; // @[bbgemm.scala 53:22]
  wire  Loop_4_clock; // @[bbgemm.scala 55:22]
  wire  Loop_4_reset; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_enable_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_enable_valid; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_enable_bits_control; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_InLiveIn_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_InLiveIn_0_valid; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_InLiveIn_0_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_InLiveIn_1_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_InLiveIn_1_valid; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_InLiveIn_1_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_InLiveIn_2_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_InLiveIn_2_valid; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_InLiveIn_2_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_activate_loop_start_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_activate_loop_start_valid; // @[bbgemm.scala 55:22]
  wire [4:0] Loop_4_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_activate_loop_start_bits_control; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_activate_loop_back_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_activate_loop_back_valid; // @[bbgemm.scala 55:22]
  wire [4:0] Loop_4_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_activate_loop_back_bits_control; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopBack_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopBack_0_valid; // @[bbgemm.scala 55:22]
  wire [4:0] Loop_4_io_loopBack_0_bits_taskID; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopBack_0_bits_control; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopFinish_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopFinish_0_valid; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopFinish_0_bits_control; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_CarryDepenIn_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_CarryDepenIn_0_valid; // @[bbgemm.scala 55:22]
  wire [4:0] Loop_4_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 55:22]
  wire [4:0] Loop_4_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 55:22]
  wire [63:0] Loop_4_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopExit_0_ready; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopExit_0_valid; // @[bbgemm.scala 55:22]
  wire [4:0] Loop_4_io_loopExit_0_bits_taskID; // @[bbgemm.scala 55:22]
  wire  Loop_4_io_loopExit_0_bits_control; // @[bbgemm.scala 55:22]
  wire  bb_entry0_clock; // @[bbgemm.scala 63:25]
  wire  bb_entry0_reset; // @[bbgemm.scala 63:25]
  wire  bb_entry0_io_predicateIn_0_ready; // @[bbgemm.scala 63:25]
  wire  bb_entry0_io_predicateIn_0_valid; // @[bbgemm.scala 63:25]
  wire  bb_entry0_io_predicateIn_0_bits_control; // @[bbgemm.scala 63:25]
  wire  bb_entry0_io_Out_0_ready; // @[bbgemm.scala 63:25]
  wire  bb_entry0_io_Out_0_valid; // @[bbgemm.scala 63:25]
  wire  bb_entry0_io_Out_0_bits_control; // @[bbgemm.scala 63:25]
  wire  bb_loopkk1_clock; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_reset; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_MaskBB_0_ready; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_MaskBB_0_valid; // @[bbgemm.scala 65:26]
  wire [1:0] bb_loopkk1_io_MaskBB_0_bits; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_0_ready; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_0_valid; // @[bbgemm.scala 65:26]
  wire [4:0] bb_loopkk1_io_Out_0_bits_taskID; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_0_bits_control; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_1_ready; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_1_valid; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_1_bits_control; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_2_ready; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_2_valid; // @[bbgemm.scala 65:26]
  wire [4:0] bb_loopkk1_io_Out_2_bits_taskID; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_Out_2_bits_control; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_predicateIn_0_ready; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_predicateIn_0_valid; // @[bbgemm.scala 65:26]
  wire [4:0] bb_loopkk1_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_predicateIn_0_bits_control; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_predicateIn_1_ready; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_predicateIn_1_valid; // @[bbgemm.scala 65:26]
  wire [4:0] bb_loopkk1_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 65:26]
  wire  bb_loopkk1_io_predicateIn_1_bits_control; // @[bbgemm.scala 65:26]
  wire  bb_loopi2_clock; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_reset; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_MaskBB_0_ready; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_MaskBB_0_valid; // @[bbgemm.scala 67:25]
  wire [1:0] bb_loopi2_io_MaskBB_0_bits; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_0_ready; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_0_valid; // @[bbgemm.scala 67:25]
  wire [4:0] bb_loopi2_io_Out_0_bits_taskID; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_0_bits_control; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_1_ready; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_1_valid; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_1_bits_control; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_2_ready; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_2_valid; // @[bbgemm.scala 67:25]
  wire [4:0] bb_loopi2_io_Out_2_bits_taskID; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_Out_2_bits_control; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_predicateIn_0_ready; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_predicateIn_0_valid; // @[bbgemm.scala 67:25]
  wire [4:0] bb_loopi2_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_predicateIn_0_bits_control; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_predicateIn_1_ready; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_predicateIn_1_valid; // @[bbgemm.scala 67:25]
  wire [4:0] bb_loopi2_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 67:25]
  wire  bb_loopi2_io_predicateIn_1_bits_control; // @[bbgemm.scala 67:25]
  wire  bb_loopk3_clock; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_reset; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_MaskBB_0_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_MaskBB_0_valid; // @[bbgemm.scala 69:25]
  wire [1:0] bb_loopk3_io_MaskBB_0_bits; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_0_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_0_valid; // @[bbgemm.scala 69:25]
  wire [4:0] bb_loopk3_io_Out_0_bits_taskID; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_0_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_1_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_1_valid; // @[bbgemm.scala 69:25]
  wire [4:0] bb_loopk3_io_Out_1_bits_taskID; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_1_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_2_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_2_valid; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_2_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_3_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_3_valid; // @[bbgemm.scala 69:25]
  wire [4:0] bb_loopk3_io_Out_3_bits_taskID; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_3_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_4_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_4_valid; // @[bbgemm.scala 69:25]
  wire [4:0] bb_loopk3_io_Out_4_bits_taskID; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_Out_4_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_predicateIn_0_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_predicateIn_0_valid; // @[bbgemm.scala 69:25]
  wire [4:0] bb_loopk3_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_predicateIn_0_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_predicateIn_1_ready; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_predicateIn_1_valid; // @[bbgemm.scala 69:25]
  wire [4:0] bb_loopk3_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 69:25]
  wire  bb_loopk3_io_predicateIn_1_bits_control; // @[bbgemm.scala 69:25]
  wire  bb_for_body94_clock; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_reset; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_MaskBB_0_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_MaskBB_0_valid; // @[bbgemm.scala 71:29]
  wire [1:0] bb_for_body94_io_MaskBB_0_bits; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_0_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_0_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_0_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_0_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_1_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_1_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_1_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_1_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_2_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_2_valid; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_2_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_3_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_3_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_3_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_3_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_4_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_4_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_4_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_4_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_5_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_5_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_5_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_5_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_6_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_6_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_6_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_6_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_7_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_7_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_7_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_7_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_8_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_8_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_8_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_8_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_9_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_9_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_Out_9_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_Out_9_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_predicateIn_0_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_predicateIn_0_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_predicateIn_0_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_predicateIn_1_ready; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_predicateIn_1_valid; // @[bbgemm.scala 71:29]
  wire [4:0] bb_for_body94_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 71:29]
  wire  bb_for_body94_io_predicateIn_1_bits_control; // @[bbgemm.scala 71:29]
  wire  bb_for_body165_clock; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_reset; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_MaskBB_0_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_MaskBB_0_valid; // @[bbgemm.scala 73:30]
  wire [1:0] bb_for_body165_io_MaskBB_0_bits; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_0_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_0_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_0_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_0_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_1_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_1_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_1_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_1_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_2_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_2_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_2_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_2_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_3_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_3_valid; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_3_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_4_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_4_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_4_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_4_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_5_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_5_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_5_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_5_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_6_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_6_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_6_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_6_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_7_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_7_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_7_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_7_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_8_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_8_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_8_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_8_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_9_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_9_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_9_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_9_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_10_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_10_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_10_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_10_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_11_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_11_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_11_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_11_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_12_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_12_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_12_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_12_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_13_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_13_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_13_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_13_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_14_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_14_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_14_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_14_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_15_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_15_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_15_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_15_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_16_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_16_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_16_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_16_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_17_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_17_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_Out_17_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_Out_17_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_predicateIn_0_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_predicateIn_0_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_predicateIn_0_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_predicateIn_1_ready; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_predicateIn_1_valid; // @[bbgemm.scala 73:30]
  wire [4:0] bb_for_body165_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 73:30]
  wire  bb_for_body165_io_predicateIn_1_bits_control; // @[bbgemm.scala 73:30]
  wire  bb_for_inc276_clock; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_reset; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_predicateIn_0_ready; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_predicateIn_0_valid; // @[bbgemm.scala 75:29]
  wire [4:0] bb_for_inc276_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_predicateIn_0_bits_control; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_0_ready; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_0_valid; // @[bbgemm.scala 75:29]
  wire [4:0] bb_for_inc276_io_Out_0_bits_taskID; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_0_bits_control; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_1_ready; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_1_valid; // @[bbgemm.scala 75:29]
  wire [4:0] bb_for_inc276_io_Out_1_bits_taskID; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_1_bits_control; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_2_ready; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_2_valid; // @[bbgemm.scala 75:29]
  wire [4:0] bb_for_inc276_io_Out_2_bits_taskID; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_2_bits_control; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_3_ready; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_3_valid; // @[bbgemm.scala 75:29]
  wire [4:0] bb_for_inc276_io_Out_3_bits_taskID; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_3_bits_control; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_4_ready; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_4_valid; // @[bbgemm.scala 75:29]
  wire [4:0] bb_for_inc276_io_Out_4_bits_taskID; // @[bbgemm.scala 75:29]
  wire  bb_for_inc276_io_Out_4_bits_control; // @[bbgemm.scala 75:29]
  wire  bb_for_inc307_clock; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_reset; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_predicateIn_0_ready; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_predicateIn_0_valid; // @[bbgemm.scala 77:29]
  wire [4:0] bb_for_inc307_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_predicateIn_0_bits_control; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_0_ready; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_0_valid; // @[bbgemm.scala 77:29]
  wire [4:0] bb_for_inc307_io_Out_0_bits_taskID; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_0_bits_control; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_1_ready; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_1_valid; // @[bbgemm.scala 77:29]
  wire [4:0] bb_for_inc307_io_Out_1_bits_taskID; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_1_bits_control; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_2_ready; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_2_valid; // @[bbgemm.scala 77:29]
  wire [4:0] bb_for_inc307_io_Out_2_bits_taskID; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_2_bits_control; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_3_ready; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_3_valid; // @[bbgemm.scala 77:29]
  wire [4:0] bb_for_inc307_io_Out_3_bits_taskID; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_3_bits_control; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_4_ready; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_4_valid; // @[bbgemm.scala 77:29]
  wire [4:0] bb_for_inc307_io_Out_4_bits_taskID; // @[bbgemm.scala 77:29]
  wire  bb_for_inc307_io_Out_4_bits_control; // @[bbgemm.scala 77:29]
  wire  bb_for_inc338_clock; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_reset; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_predicateIn_0_ready; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_predicateIn_0_valid; // @[bbgemm.scala 79:29]
  wire [4:0] bb_for_inc338_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_predicateIn_0_bits_control; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_0_ready; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_0_valid; // @[bbgemm.scala 79:29]
  wire [4:0] bb_for_inc338_io_Out_0_bits_taskID; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_0_bits_control; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_1_ready; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_1_valid; // @[bbgemm.scala 79:29]
  wire [4:0] bb_for_inc338_io_Out_1_bits_taskID; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_1_bits_control; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_2_ready; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_2_valid; // @[bbgemm.scala 79:29]
  wire [4:0] bb_for_inc338_io_Out_2_bits_taskID; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_2_bits_control; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_3_ready; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_3_valid; // @[bbgemm.scala 79:29]
  wire [4:0] bb_for_inc338_io_Out_3_bits_taskID; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_3_bits_control; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_4_ready; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_4_valid; // @[bbgemm.scala 79:29]
  wire [4:0] bb_for_inc338_io_Out_4_bits_taskID; // @[bbgemm.scala 79:29]
  wire  bb_for_inc338_io_Out_4_bits_control; // @[bbgemm.scala 79:29]
  wire  bb_for_inc369_clock; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_reset; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_predicateIn_0_ready; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_predicateIn_0_valid; // @[bbgemm.scala 81:29]
  wire [4:0] bb_for_inc369_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_predicateIn_0_bits_control; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_0_ready; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_0_valid; // @[bbgemm.scala 81:29]
  wire [4:0] bb_for_inc369_io_Out_0_bits_taskID; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_0_bits_control; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_1_ready; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_1_valid; // @[bbgemm.scala 81:29]
  wire [4:0] bb_for_inc369_io_Out_1_bits_taskID; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_1_bits_control; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_2_ready; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_2_valid; // @[bbgemm.scala 81:29]
  wire [4:0] bb_for_inc369_io_Out_2_bits_taskID; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_2_bits_control; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_3_ready; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_3_valid; // @[bbgemm.scala 81:29]
  wire [4:0] bb_for_inc369_io_Out_3_bits_taskID; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_3_bits_control; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_4_ready; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_4_valid; // @[bbgemm.scala 81:29]
  wire [4:0] bb_for_inc369_io_Out_4_bits_taskID; // @[bbgemm.scala 81:29]
  wire  bb_for_inc369_io_Out_4_bits_control; // @[bbgemm.scala 81:29]
  wire  bb_for_end3810_clock; // @[bbgemm.scala 83:30]
  wire  bb_for_end3810_reset; // @[bbgemm.scala 83:30]
  wire  bb_for_end3810_io_predicateIn_0_ready; // @[bbgemm.scala 83:30]
  wire  bb_for_end3810_io_predicateIn_0_valid; // @[bbgemm.scala 83:30]
  wire [4:0] bb_for_end3810_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 83:30]
  wire  bb_for_end3810_io_predicateIn_0_bits_control; // @[bbgemm.scala 83:30]
  wire  bb_for_end3810_io_Out_0_ready; // @[bbgemm.scala 83:30]
  wire  bb_for_end3810_io_Out_0_valid; // @[bbgemm.scala 83:30]
  wire [4:0] bb_for_end3810_io_Out_0_bits_taskID; // @[bbgemm.scala 83:30]
  wire  br_0_clock; // @[bbgemm.scala 92:20]
  wire  br_0_reset; // @[bbgemm.scala 92:20]
  wire  br_0_io_enable_ready; // @[bbgemm.scala 92:20]
  wire  br_0_io_enable_valid; // @[bbgemm.scala 92:20]
  wire  br_0_io_enable_bits_control; // @[bbgemm.scala 92:20]
  wire  br_0_io_Out_0_ready; // @[bbgemm.scala 92:20]
  wire  br_0_io_Out_0_valid; // @[bbgemm.scala 92:20]
  wire  br_0_io_Out_0_bits_control; // @[bbgemm.scala 92:20]
  wire  phiindvars_iv841_clock; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_reset; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_enable_ready; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_enable_valid; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_enable_bits_control; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_InData_0_ready; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_InData_0_valid; // @[bbgemm.scala 95:32]
  wire [4:0] phiindvars_iv841_io_InData_0_bits_taskID; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_InData_1_ready; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_InData_1_valid; // @[bbgemm.scala 95:32]
  wire [4:0] phiindvars_iv841_io_InData_1_bits_taskID; // @[bbgemm.scala 95:32]
  wire [63:0] phiindvars_iv841_io_InData_1_bits_data; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_Mask_ready; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_Mask_valid; // @[bbgemm.scala 95:32]
  wire [1:0] phiindvars_iv841_io_Mask_bits; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_Out_0_ready; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_Out_0_valid; // @[bbgemm.scala 95:32]
  wire [63:0] phiindvars_iv841_io_Out_0_bits_data; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_Out_1_ready; // @[bbgemm.scala 95:32]
  wire  phiindvars_iv841_io_Out_1_valid; // @[bbgemm.scala 95:32]
  wire [63:0] phiindvars_iv841_io_Out_1_bits_data; // @[bbgemm.scala 95:32]
  wire  br_2_clock; // @[bbgemm.scala 97:20]
  wire  br_2_reset; // @[bbgemm.scala 97:20]
  wire  br_2_io_enable_ready; // @[bbgemm.scala 97:20]
  wire  br_2_io_enable_valid; // @[bbgemm.scala 97:20]
  wire [4:0] br_2_io_enable_bits_taskID; // @[bbgemm.scala 97:20]
  wire  br_2_io_enable_bits_control; // @[bbgemm.scala 97:20]
  wire  br_2_io_Out_0_ready; // @[bbgemm.scala 97:20]
  wire  br_2_io_Out_0_valid; // @[bbgemm.scala 97:20]
  wire [4:0] br_2_io_Out_0_bits_taskID; // @[bbgemm.scala 97:20]
  wire  br_2_io_Out_0_bits_control; // @[bbgemm.scala 97:20]
  wire  phiindvars_iv823_clock; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_reset; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_enable_ready; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_enable_valid; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_enable_bits_control; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_InData_0_ready; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_InData_0_valid; // @[bbgemm.scala 100:32]
  wire [4:0] phiindvars_iv823_io_InData_0_bits_taskID; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_InData_1_ready; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_InData_1_valid; // @[bbgemm.scala 100:32]
  wire [4:0] phiindvars_iv823_io_InData_1_bits_taskID; // @[bbgemm.scala 100:32]
  wire [63:0] phiindvars_iv823_io_InData_1_bits_data; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_Mask_ready; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_Mask_valid; // @[bbgemm.scala 100:32]
  wire [1:0] phiindvars_iv823_io_Mask_bits; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_Out_0_ready; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_Out_0_valid; // @[bbgemm.scala 100:32]
  wire [63:0] phiindvars_iv823_io_Out_0_bits_data; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_Out_1_ready; // @[bbgemm.scala 100:32]
  wire  phiindvars_iv823_io_Out_1_valid; // @[bbgemm.scala 100:32]
  wire [63:0] phiindvars_iv823_io_Out_1_bits_data; // @[bbgemm.scala 100:32]
  wire  br_4_clock; // @[bbgemm.scala 104:20]
  wire  br_4_reset; // @[bbgemm.scala 104:20]
  wire  br_4_io_enable_ready; // @[bbgemm.scala 104:20]
  wire  br_4_io_enable_valid; // @[bbgemm.scala 104:20]
  wire [4:0] br_4_io_enable_bits_taskID; // @[bbgemm.scala 104:20]
  wire  br_4_io_enable_bits_control; // @[bbgemm.scala 104:20]
  wire  br_4_io_Out_0_ready; // @[bbgemm.scala 104:20]
  wire  br_4_io_Out_0_valid; // @[bbgemm.scala 104:20]
  wire [4:0] br_4_io_Out_0_bits_taskID; // @[bbgemm.scala 104:20]
  wire  br_4_io_Out_0_bits_control; // @[bbgemm.scala 104:20]
  wire  phiindvars_iv785_clock; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_reset; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_enable_ready; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_enable_valid; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_enable_bits_control; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_InData_0_ready; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_InData_0_valid; // @[bbgemm.scala 107:32]
  wire [4:0] phiindvars_iv785_io_InData_0_bits_taskID; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_InData_1_ready; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_InData_1_valid; // @[bbgemm.scala 107:32]
  wire [4:0] phiindvars_iv785_io_InData_1_bits_taskID; // @[bbgemm.scala 107:32]
  wire [63:0] phiindvars_iv785_io_InData_1_bits_data; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_Mask_ready; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_Mask_valid; // @[bbgemm.scala 107:32]
  wire [1:0] phiindvars_iv785_io_Mask_bits; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_Out_0_ready; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_Out_0_valid; // @[bbgemm.scala 107:32]
  wire [63:0] phiindvars_iv785_io_Out_0_bits_data; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_Out_1_ready; // @[bbgemm.scala 107:32]
  wire  phiindvars_iv785_io_Out_1_valid; // @[bbgemm.scala 107:32]
  wire [63:0] phiindvars_iv785_io_Out_1_bits_data; // @[bbgemm.scala 107:32]
  wire  binaryOp_6_clock; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_reset; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_enable_ready; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_enable_valid; // @[bbgemm.scala 119:26]
  wire [4:0] binaryOp_6_io_enable_bits_taskID; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_enable_bits_control; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_Out_0_ready; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_Out_0_valid; // @[bbgemm.scala 119:26]
  wire [63:0] binaryOp_6_io_Out_0_bits_data; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_LeftIO_ready; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_LeftIO_valid; // @[bbgemm.scala 119:26]
  wire [63:0] binaryOp_6_io_LeftIO_bits_data; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_RightIO_ready; // @[bbgemm.scala 119:26]
  wire  binaryOp_6_io_RightIO_valid; // @[bbgemm.scala 119:26]
  wire  br_7_clock; // @[bbgemm.scala 122:20]
  wire  br_7_reset; // @[bbgemm.scala 122:20]
  wire  br_7_io_enable_ready; // @[bbgemm.scala 122:20]
  wire  br_7_io_enable_valid; // @[bbgemm.scala 122:20]
  wire [4:0] br_7_io_enable_bits_taskID; // @[bbgemm.scala 122:20]
  wire  br_7_io_enable_bits_control; // @[bbgemm.scala 122:20]
  wire  br_7_io_Out_0_ready; // @[bbgemm.scala 122:20]
  wire  br_7_io_Out_0_valid; // @[bbgemm.scala 122:20]
  wire [4:0] br_7_io_Out_0_bits_taskID; // @[bbgemm.scala 122:20]
  wire  br_7_io_Out_0_bits_control; // @[bbgemm.scala 122:20]
  wire  phiindvars_iv718_clock; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_reset; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_enable_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_enable_valid; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_enable_bits_control; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_InData_0_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_InData_0_valid; // @[bbgemm.scala 125:32]
  wire [4:0] phiindvars_iv718_io_InData_0_bits_taskID; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_InData_1_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_InData_1_valid; // @[bbgemm.scala 125:32]
  wire [4:0] phiindvars_iv718_io_InData_1_bits_taskID; // @[bbgemm.scala 125:32]
  wire [63:0] phiindvars_iv718_io_InData_1_bits_data; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Mask_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Mask_valid; // @[bbgemm.scala 125:32]
  wire [1:0] phiindvars_iv718_io_Mask_bits; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Out_0_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Out_0_valid; // @[bbgemm.scala 125:32]
  wire [63:0] phiindvars_iv718_io_Out_0_bits_data; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Out_1_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Out_1_valid; // @[bbgemm.scala 125:32]
  wire [63:0] phiindvars_iv718_io_Out_1_bits_data; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Out_2_ready; // @[bbgemm.scala 125:32]
  wire  phiindvars_iv718_io_Out_2_valid; // @[bbgemm.scala 125:32]
  wire [63:0] phiindvars_iv718_io_Out_2_bits_data; // @[bbgemm.scala 125:32]
  wire  binaryOp_9_clock; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_reset; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_enable_ready; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_enable_valid; // @[bbgemm.scala 128:26]
  wire [4:0] binaryOp_9_io_enable_bits_taskID; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_enable_bits_control; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_Out_0_ready; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_Out_0_valid; // @[bbgemm.scala 128:26]
  wire [63:0] binaryOp_9_io_Out_0_bits_data; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_LeftIO_ready; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_LeftIO_valid; // @[bbgemm.scala 128:26]
  wire [63:0] binaryOp_9_io_LeftIO_bits_data; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_RightIO_ready; // @[bbgemm.scala 128:26]
  wire  binaryOp_9_io_RightIO_valid; // @[bbgemm.scala 128:26]
  wire [63:0] binaryOp_9_io_RightIO_bits_data; // @[bbgemm.scala 128:26]
  wire  binaryOp_10_clock; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_reset; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_enable_ready; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_enable_valid; // @[bbgemm.scala 131:27]
  wire [4:0] binaryOp_10_io_enable_bits_taskID; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_enable_bits_control; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_Out_0_ready; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_Out_0_valid; // @[bbgemm.scala 131:27]
  wire [63:0] binaryOp_10_io_Out_0_bits_data; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_LeftIO_ready; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_LeftIO_valid; // @[bbgemm.scala 131:27]
  wire [63:0] binaryOp_10_io_LeftIO_bits_data; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_RightIO_ready; // @[bbgemm.scala 131:27]
  wire  binaryOp_10_io_RightIO_valid; // @[bbgemm.scala 131:27]
  wire  binaryOp_11_clock; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_reset; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_enable_ready; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_enable_valid; // @[bbgemm.scala 134:27]
  wire [4:0] binaryOp_11_io_enable_bits_taskID; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_enable_bits_control; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_Out_0_ready; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_Out_0_valid; // @[bbgemm.scala 134:27]
  wire [63:0] binaryOp_11_io_Out_0_bits_data; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_LeftIO_ready; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_LeftIO_valid; // @[bbgemm.scala 134:27]
  wire [63:0] binaryOp_11_io_LeftIO_bits_data; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_RightIO_ready; // @[bbgemm.scala 134:27]
  wire  binaryOp_11_io_RightIO_valid; // @[bbgemm.scala 134:27]
  wire [63:0] binaryOp_11_io_RightIO_bits_data; // @[bbgemm.scala 134:27]
  wire  binaryOp_12_clock; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_reset; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_enable_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_enable_valid; // @[bbgemm.scala 137:27]
  wire [4:0] binaryOp_12_io_enable_bits_taskID; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_enable_bits_control; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_Out_0_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_Out_0_valid; // @[bbgemm.scala 137:27]
  wire [63:0] binaryOp_12_io_Out_0_bits_data; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_LeftIO_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_LeftIO_valid; // @[bbgemm.scala 137:27]
  wire [63:0] binaryOp_12_io_LeftIO_bits_data; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_RightIO_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_12_io_RightIO_valid; // @[bbgemm.scala 137:27]
  wire [63:0] binaryOp_12_io_RightIO_bits_data; // @[bbgemm.scala 137:27]
  wire  Gep_arrayidx13_clock; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_reset; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_enable_ready; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_enable_valid; // @[bbgemm.scala 140:30]
  wire [4:0] Gep_arrayidx13_io_enable_bits_taskID; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_enable_bits_control; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_Out_0_ready; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_Out_0_valid; // @[bbgemm.scala 140:30]
  wire [63:0] Gep_arrayidx13_io_Out_0_bits_data; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_baseAddress_ready; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_baseAddress_valid; // @[bbgemm.scala 140:30]
  wire [63:0] Gep_arrayidx13_io_baseAddress_bits_data; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_idx_0_ready; // @[bbgemm.scala 140:30]
  wire  Gep_arrayidx13_io_idx_0_valid; // @[bbgemm.scala 140:30]
  wire [63:0] Gep_arrayidx13_io_idx_0_bits_data; // @[bbgemm.scala 140:30]
  wire  ld_14_clock; // @[bbgemm.scala 143:21]
  wire  ld_14_reset; // @[bbgemm.scala 143:21]
  wire  ld_14_io_enable_ready; // @[bbgemm.scala 143:21]
  wire  ld_14_io_enable_valid; // @[bbgemm.scala 143:21]
  wire [4:0] ld_14_io_enable_bits_taskID; // @[bbgemm.scala 143:21]
  wire  ld_14_io_enable_bits_control; // @[bbgemm.scala 143:21]
  wire  ld_14_io_Out_0_ready; // @[bbgemm.scala 143:21]
  wire  ld_14_io_Out_0_valid; // @[bbgemm.scala 143:21]
  wire [63:0] ld_14_io_Out_0_bits_data; // @[bbgemm.scala 143:21]
  wire  ld_14_io_GepAddr_ready; // @[bbgemm.scala 143:21]
  wire  ld_14_io_GepAddr_valid; // @[bbgemm.scala 143:21]
  wire [63:0] ld_14_io_GepAddr_bits_data; // @[bbgemm.scala 143:21]
  wire  ld_14_io_MemReq_ready; // @[bbgemm.scala 143:21]
  wire  ld_14_io_MemReq_valid; // @[bbgemm.scala 143:21]
  wire [63:0] ld_14_io_MemReq_bits_addr; // @[bbgemm.scala 143:21]
  wire  ld_14_io_MemResp_valid; // @[bbgemm.scala 143:21]
  wire [63:0] ld_14_io_MemResp_bits_data; // @[bbgemm.scala 143:21]
  wire  br_15_clock; // @[bbgemm.scala 146:21]
  wire  br_15_reset; // @[bbgemm.scala 146:21]
  wire  br_15_io_enable_ready; // @[bbgemm.scala 146:21]
  wire  br_15_io_enable_valid; // @[bbgemm.scala 146:21]
  wire [4:0] br_15_io_enable_bits_taskID; // @[bbgemm.scala 146:21]
  wire  br_15_io_enable_bits_control; // @[bbgemm.scala 146:21]
  wire  br_15_io_Out_0_ready; // @[bbgemm.scala 146:21]
  wire  br_15_io_Out_0_valid; // @[bbgemm.scala 146:21]
  wire [4:0] br_15_io_Out_0_bits_taskID; // @[bbgemm.scala 146:21]
  wire  br_15_io_Out_0_bits_control; // @[bbgemm.scala 146:21]
  wire  phiindvars_iv16_clock; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_reset; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_enable_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_enable_valid; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_enable_bits_control; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_InData_0_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_InData_0_valid; // @[bbgemm.scala 149:31]
  wire [4:0] phiindvars_iv16_io_InData_0_bits_taskID; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_InData_1_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_InData_1_valid; // @[bbgemm.scala 149:31]
  wire [4:0] phiindvars_iv16_io_InData_1_bits_taskID; // @[bbgemm.scala 149:31]
  wire [63:0] phiindvars_iv16_io_InData_1_bits_data; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Mask_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Mask_valid; // @[bbgemm.scala 149:31]
  wire [1:0] phiindvars_iv16_io_Mask_bits; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Out_0_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Out_0_valid; // @[bbgemm.scala 149:31]
  wire [63:0] phiindvars_iv16_io_Out_0_bits_data; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Out_1_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Out_1_valid; // @[bbgemm.scala 149:31]
  wire [63:0] phiindvars_iv16_io_Out_1_bits_data; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Out_2_ready; // @[bbgemm.scala 149:31]
  wire  phiindvars_iv16_io_Out_2_valid; // @[bbgemm.scala 149:31]
  wire [63:0] phiindvars_iv16_io_Out_2_bits_data; // @[bbgemm.scala 149:31]
  wire  binaryOp_17_clock; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_reset; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_enable_ready; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_enable_valid; // @[bbgemm.scala 152:27]
  wire [4:0] binaryOp_17_io_enable_bits_taskID; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_enable_bits_control; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_Out_0_ready; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_Out_0_valid; // @[bbgemm.scala 152:27]
  wire [63:0] binaryOp_17_io_Out_0_bits_data; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_LeftIO_ready; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_LeftIO_valid; // @[bbgemm.scala 152:27]
  wire [63:0] binaryOp_17_io_LeftIO_bits_data; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_RightIO_ready; // @[bbgemm.scala 152:27]
  wire  binaryOp_17_io_RightIO_valid; // @[bbgemm.scala 152:27]
  wire [63:0] binaryOp_17_io_RightIO_bits_data; // @[bbgemm.scala 152:27]
  wire  binaryOp_18_clock; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_reset; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_enable_ready; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_enable_valid; // @[bbgemm.scala 155:27]
  wire [4:0] binaryOp_18_io_enable_bits_taskID; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_enable_bits_control; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_Out_0_ready; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_Out_0_valid; // @[bbgemm.scala 155:27]
  wire [63:0] binaryOp_18_io_Out_0_bits_data; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_LeftIO_ready; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_LeftIO_valid; // @[bbgemm.scala 155:27]
  wire [63:0] binaryOp_18_io_LeftIO_bits_data; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_RightIO_ready; // @[bbgemm.scala 155:27]
  wire  binaryOp_18_io_RightIO_valid; // @[bbgemm.scala 155:27]
  wire [63:0] binaryOp_18_io_RightIO_bits_data; // @[bbgemm.scala 155:27]
  wire  Gep_arrayidx2019_clock; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_reset; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_enable_ready; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_enable_valid; // @[bbgemm.scala 158:32]
  wire [4:0] Gep_arrayidx2019_io_enable_bits_taskID; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_enable_bits_control; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_Out_0_ready; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_Out_0_valid; // @[bbgemm.scala 158:32]
  wire [63:0] Gep_arrayidx2019_io_Out_0_bits_data; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_baseAddress_ready; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_baseAddress_valid; // @[bbgemm.scala 158:32]
  wire [63:0] Gep_arrayidx2019_io_baseAddress_bits_data; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_idx_0_ready; // @[bbgemm.scala 158:32]
  wire  Gep_arrayidx2019_io_idx_0_valid; // @[bbgemm.scala 158:32]
  wire [63:0] Gep_arrayidx2019_io_idx_0_bits_data; // @[bbgemm.scala 158:32]
  wire  ld_20_clock; // @[bbgemm.scala 161:21]
  wire  ld_20_reset; // @[bbgemm.scala 161:21]
  wire  ld_20_io_enable_ready; // @[bbgemm.scala 161:21]
  wire  ld_20_io_enable_valid; // @[bbgemm.scala 161:21]
  wire [4:0] ld_20_io_enable_bits_taskID; // @[bbgemm.scala 161:21]
  wire  ld_20_io_enable_bits_control; // @[bbgemm.scala 161:21]
  wire  ld_20_io_Out_0_ready; // @[bbgemm.scala 161:21]
  wire  ld_20_io_Out_0_valid; // @[bbgemm.scala 161:21]
  wire [63:0] ld_20_io_Out_0_bits_data; // @[bbgemm.scala 161:21]
  wire  ld_20_io_GepAddr_ready; // @[bbgemm.scala 161:21]
  wire  ld_20_io_GepAddr_valid; // @[bbgemm.scala 161:21]
  wire [63:0] ld_20_io_GepAddr_bits_data; // @[bbgemm.scala 161:21]
  wire  ld_20_io_MemReq_ready; // @[bbgemm.scala 161:21]
  wire  ld_20_io_MemReq_valid; // @[bbgemm.scala 161:21]
  wire [63:0] ld_20_io_MemReq_bits_addr; // @[bbgemm.scala 161:21]
  wire  ld_20_io_MemResp_valid; // @[bbgemm.scala 161:21]
  wire [63:0] ld_20_io_MemResp_bits_data; // @[bbgemm.scala 161:21]
  wire  FP_mul2121_clock; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_reset; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_enable_ready; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_enable_valid; // @[bbgemm.scala 164:26]
  wire [4:0] FP_mul2121_io_enable_bits_taskID; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_enable_bits_control; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_Out_0_ready; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_Out_0_valid; // @[bbgemm.scala 164:26]
  wire [63:0] FP_mul2121_io_Out_0_bits_data; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_LeftIO_ready; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_LeftIO_valid; // @[bbgemm.scala 164:26]
  wire [63:0] FP_mul2121_io_LeftIO_bits_data; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_RightIO_ready; // @[bbgemm.scala 164:26]
  wire  FP_mul2121_io_RightIO_valid; // @[bbgemm.scala 164:26]
  wire [63:0] FP_mul2121_io_RightIO_bits_data; // @[bbgemm.scala 164:26]
  wire  binaryOp_22_clock; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_reset; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_enable_ready; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_enable_valid; // @[bbgemm.scala 167:27]
  wire [4:0] binaryOp_22_io_enable_bits_taskID; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_enable_bits_control; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_Out_0_ready; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_Out_0_valid; // @[bbgemm.scala 167:27]
  wire [63:0] binaryOp_22_io_Out_0_bits_data; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_LeftIO_ready; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_LeftIO_valid; // @[bbgemm.scala 167:27]
  wire [63:0] binaryOp_22_io_LeftIO_bits_data; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_RightIO_ready; // @[bbgemm.scala 167:27]
  wire  binaryOp_22_io_RightIO_valid; // @[bbgemm.scala 167:27]
  wire [63:0] binaryOp_22_io_RightIO_bits_data; // @[bbgemm.scala 167:27]
  wire  binaryOp_23_clock; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_reset; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_enable_ready; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_enable_valid; // @[bbgemm.scala 170:27]
  wire [4:0] binaryOp_23_io_enable_bits_taskID; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_enable_bits_control; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_Out_0_ready; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_Out_0_valid; // @[bbgemm.scala 170:27]
  wire [63:0] binaryOp_23_io_Out_0_bits_data; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_LeftIO_ready; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_LeftIO_valid; // @[bbgemm.scala 170:27]
  wire [63:0] binaryOp_23_io_LeftIO_bits_data; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_RightIO_ready; // @[bbgemm.scala 170:27]
  wire  binaryOp_23_io_RightIO_valid; // @[bbgemm.scala 170:27]
  wire [63:0] binaryOp_23_io_RightIO_bits_data; // @[bbgemm.scala 170:27]
  wire  Gep_arrayidx2524_clock; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_reset; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_enable_ready; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_enable_valid; // @[bbgemm.scala 173:32]
  wire [4:0] Gep_arrayidx2524_io_enable_bits_taskID; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_enable_bits_control; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_Out_0_ready; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_Out_0_valid; // @[bbgemm.scala 173:32]
  wire [63:0] Gep_arrayidx2524_io_Out_0_bits_data; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_Out_1_ready; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_Out_1_valid; // @[bbgemm.scala 173:32]
  wire [63:0] Gep_arrayidx2524_io_Out_1_bits_data; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_baseAddress_ready; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_baseAddress_valid; // @[bbgemm.scala 173:32]
  wire [63:0] Gep_arrayidx2524_io_baseAddress_bits_data; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_idx_0_ready; // @[bbgemm.scala 173:32]
  wire  Gep_arrayidx2524_io_idx_0_valid; // @[bbgemm.scala 173:32]
  wire [63:0] Gep_arrayidx2524_io_idx_0_bits_data; // @[bbgemm.scala 173:32]
  wire  ld_25_clock; // @[bbgemm.scala 176:21]
  wire  ld_25_reset; // @[bbgemm.scala 176:21]
  wire  ld_25_io_enable_ready; // @[bbgemm.scala 176:21]
  wire  ld_25_io_enable_valid; // @[bbgemm.scala 176:21]
  wire [4:0] ld_25_io_enable_bits_taskID; // @[bbgemm.scala 176:21]
  wire  ld_25_io_enable_bits_control; // @[bbgemm.scala 176:21]
  wire  ld_25_io_Out_0_ready; // @[bbgemm.scala 176:21]
  wire  ld_25_io_Out_0_valid; // @[bbgemm.scala 176:21]
  wire [63:0] ld_25_io_Out_0_bits_data; // @[bbgemm.scala 176:21]
  wire  ld_25_io_GepAddr_ready; // @[bbgemm.scala 176:21]
  wire  ld_25_io_GepAddr_valid; // @[bbgemm.scala 176:21]
  wire [63:0] ld_25_io_GepAddr_bits_data; // @[bbgemm.scala 176:21]
  wire  ld_25_io_MemReq_ready; // @[bbgemm.scala 176:21]
  wire  ld_25_io_MemReq_valid; // @[bbgemm.scala 176:21]
  wire [63:0] ld_25_io_MemReq_bits_addr; // @[bbgemm.scala 176:21]
  wire  ld_25_io_MemResp_valid; // @[bbgemm.scala 176:21]
  wire [63:0] ld_25_io_MemResp_bits_data; // @[bbgemm.scala 176:21]
  wire  FP_add2626_clock; // @[bbgemm.scala 179:26]
  wire  FP_add2626_reset; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_enable_ready; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_enable_valid; // @[bbgemm.scala 179:26]
  wire [4:0] FP_add2626_io_enable_bits_taskID; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_enable_bits_control; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_Out_0_ready; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_Out_0_valid; // @[bbgemm.scala 179:26]
  wire [63:0] FP_add2626_io_Out_0_bits_data; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_LeftIO_ready; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_LeftIO_valid; // @[bbgemm.scala 179:26]
  wire [63:0] FP_add2626_io_LeftIO_bits_data; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_RightIO_ready; // @[bbgemm.scala 179:26]
  wire  FP_add2626_io_RightIO_valid; // @[bbgemm.scala 179:26]
  wire [63:0] FP_add2626_io_RightIO_bits_data; // @[bbgemm.scala 179:26]
  wire  st_27_clock; // @[bbgemm.scala 182:21]
  wire  st_27_reset; // @[bbgemm.scala 182:21]
  wire  st_27_io_enable_ready; // @[bbgemm.scala 182:21]
  wire  st_27_io_enable_valid; // @[bbgemm.scala 182:21]
  wire [4:0] st_27_io_enable_bits_taskID; // @[bbgemm.scala 182:21]
  wire  st_27_io_enable_bits_control; // @[bbgemm.scala 182:21]
  wire  st_27_io_SuccOp_0_ready; // @[bbgemm.scala 182:21]
  wire  st_27_io_SuccOp_0_valid; // @[bbgemm.scala 182:21]
  wire  st_27_io_GepAddr_ready; // @[bbgemm.scala 182:21]
  wire  st_27_io_GepAddr_valid; // @[bbgemm.scala 182:21]
  wire [63:0] st_27_io_GepAddr_bits_data; // @[bbgemm.scala 182:21]
  wire  st_27_io_inData_ready; // @[bbgemm.scala 182:21]
  wire  st_27_io_inData_valid; // @[bbgemm.scala 182:21]
  wire [63:0] st_27_io_inData_bits_data; // @[bbgemm.scala 182:21]
  wire  st_27_io_MemReq_ready; // @[bbgemm.scala 182:21]
  wire  st_27_io_MemReq_valid; // @[bbgemm.scala 182:21]
  wire [63:0] st_27_io_MemReq_bits_addr; // @[bbgemm.scala 182:21]
  wire [63:0] st_27_io_MemReq_bits_data; // @[bbgemm.scala 182:21]
  wire  st_27_io_MemResp_valid; // @[bbgemm.scala 182:21]
  wire  binaryOp_indvars_iv_next28_clock; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_reset; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_enable_ready; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_enable_valid; // @[bbgemm.scala 185:42]
  wire [4:0] binaryOp_indvars_iv_next28_io_enable_bits_taskID; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_enable_bits_control; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_Out_0_ready; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_Out_0_valid; // @[bbgemm.scala 185:42]
  wire [4:0] binaryOp_indvars_iv_next28_io_Out_0_bits_taskID; // @[bbgemm.scala 185:42]
  wire [63:0] binaryOp_indvars_iv_next28_io_Out_0_bits_data; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_Out_1_ready; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_Out_1_valid; // @[bbgemm.scala 185:42]
  wire [63:0] binaryOp_indvars_iv_next28_io_Out_1_bits_data; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_LeftIO_ready; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_LeftIO_valid; // @[bbgemm.scala 185:42]
  wire [63:0] binaryOp_indvars_iv_next28_io_LeftIO_bits_data; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_RightIO_ready; // @[bbgemm.scala 185:42]
  wire  binaryOp_indvars_iv_next28_io_RightIO_valid; // @[bbgemm.scala 185:42]
  wire  icmp_exitcond29_clock; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_reset; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_enable_ready; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_enable_valid; // @[bbgemm.scala 188:31]
  wire [4:0] icmp_exitcond29_io_enable_bits_taskID; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_enable_bits_control; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_Out_0_ready; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_Out_0_valid; // @[bbgemm.scala 188:31]
  wire [4:0] icmp_exitcond29_io_Out_0_bits_taskID; // @[bbgemm.scala 188:31]
  wire [63:0] icmp_exitcond29_io_Out_0_bits_data; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_LeftIO_ready; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_LeftIO_valid; // @[bbgemm.scala 188:31]
  wire [63:0] icmp_exitcond29_io_LeftIO_bits_data; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_RightIO_ready; // @[bbgemm.scala 188:31]
  wire  icmp_exitcond29_io_RightIO_valid; // @[bbgemm.scala 188:31]
  wire  br_30_clock; // @[bbgemm.scala 191:21]
  wire  br_30_reset; // @[bbgemm.scala 191:21]
  wire  br_30_io_enable_ready; // @[bbgemm.scala 191:21]
  wire  br_30_io_enable_valid; // @[bbgemm.scala 191:21]
  wire [4:0] br_30_io_enable_bits_taskID; // @[bbgemm.scala 191:21]
  wire  br_30_io_enable_bits_control; // @[bbgemm.scala 191:21]
  wire  br_30_io_CmpIO_ready; // @[bbgemm.scala 191:21]
  wire  br_30_io_CmpIO_valid; // @[bbgemm.scala 191:21]
  wire [4:0] br_30_io_CmpIO_bits_taskID; // @[bbgemm.scala 191:21]
  wire [63:0] br_30_io_CmpIO_bits_data; // @[bbgemm.scala 191:21]
  wire  br_30_io_PredOp_0_ready; // @[bbgemm.scala 191:21]
  wire  br_30_io_PredOp_0_valid; // @[bbgemm.scala 191:21]
  wire  br_30_io_TrueOutput_0_ready; // @[bbgemm.scala 191:21]
  wire  br_30_io_TrueOutput_0_valid; // @[bbgemm.scala 191:21]
  wire  br_30_io_TrueOutput_0_bits_control; // @[bbgemm.scala 191:21]
  wire  br_30_io_FalseOutput_0_ready; // @[bbgemm.scala 191:21]
  wire  br_30_io_FalseOutput_0_valid; // @[bbgemm.scala 191:21]
  wire [4:0] br_30_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 191:21]
  wire  br_30_io_FalseOutput_0_bits_control; // @[bbgemm.scala 191:21]
  wire  binaryOp_indvars_iv_next7231_clock; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_reset; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_enable_ready; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_enable_valid; // @[bbgemm.scala 194:44]
  wire [4:0] binaryOp_indvars_iv_next7231_io_enable_bits_taskID; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_enable_bits_control; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_Out_0_ready; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_Out_0_valid; // @[bbgemm.scala 194:44]
  wire [4:0] binaryOp_indvars_iv_next7231_io_Out_0_bits_taskID; // @[bbgemm.scala 194:44]
  wire [63:0] binaryOp_indvars_iv_next7231_io_Out_0_bits_data; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_Out_1_ready; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_Out_1_valid; // @[bbgemm.scala 194:44]
  wire [63:0] binaryOp_indvars_iv_next7231_io_Out_1_bits_data; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_LeftIO_ready; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_LeftIO_valid; // @[bbgemm.scala 194:44]
  wire [63:0] binaryOp_indvars_iv_next7231_io_LeftIO_bits_data; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_RightIO_ready; // @[bbgemm.scala 194:44]
  wire  binaryOp_indvars_iv_next7231_io_RightIO_valid; // @[bbgemm.scala 194:44]
  wire  icmp_exitcond7732_clock; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_reset; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_enable_ready; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_enable_valid; // @[bbgemm.scala 197:33]
  wire [4:0] icmp_exitcond7732_io_enable_bits_taskID; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_enable_bits_control; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_Out_0_ready; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_Out_0_valid; // @[bbgemm.scala 197:33]
  wire [4:0] icmp_exitcond7732_io_Out_0_bits_taskID; // @[bbgemm.scala 197:33]
  wire [63:0] icmp_exitcond7732_io_Out_0_bits_data; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_LeftIO_ready; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_LeftIO_valid; // @[bbgemm.scala 197:33]
  wire [63:0] icmp_exitcond7732_io_LeftIO_bits_data; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_RightIO_ready; // @[bbgemm.scala 197:33]
  wire  icmp_exitcond7732_io_RightIO_valid; // @[bbgemm.scala 197:33]
  wire  br_33_clock; // @[bbgemm.scala 200:21]
  wire  br_33_reset; // @[bbgemm.scala 200:21]
  wire  br_33_io_enable_ready; // @[bbgemm.scala 200:21]
  wire  br_33_io_enable_valid; // @[bbgemm.scala 200:21]
  wire [4:0] br_33_io_enable_bits_taskID; // @[bbgemm.scala 200:21]
  wire  br_33_io_enable_bits_control; // @[bbgemm.scala 200:21]
  wire  br_33_io_CmpIO_ready; // @[bbgemm.scala 200:21]
  wire  br_33_io_CmpIO_valid; // @[bbgemm.scala 200:21]
  wire [4:0] br_33_io_CmpIO_bits_taskID; // @[bbgemm.scala 200:21]
  wire [63:0] br_33_io_CmpIO_bits_data; // @[bbgemm.scala 200:21]
  wire  br_33_io_TrueOutput_0_ready; // @[bbgemm.scala 200:21]
  wire  br_33_io_TrueOutput_0_valid; // @[bbgemm.scala 200:21]
  wire  br_33_io_TrueOutput_0_bits_control; // @[bbgemm.scala 200:21]
  wire  br_33_io_FalseOutput_0_ready; // @[bbgemm.scala 200:21]
  wire  br_33_io_FalseOutput_0_valid; // @[bbgemm.scala 200:21]
  wire [4:0] br_33_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 200:21]
  wire  br_33_io_FalseOutput_0_bits_control; // @[bbgemm.scala 200:21]
  wire  binaryOp_indvars_iv_next7934_clock; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_reset; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_enable_ready; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_enable_valid; // @[bbgemm.scala 203:44]
  wire [4:0] binaryOp_indvars_iv_next7934_io_enable_bits_taskID; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_enable_bits_control; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_Out_0_ready; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_Out_0_valid; // @[bbgemm.scala 203:44]
  wire [4:0] binaryOp_indvars_iv_next7934_io_Out_0_bits_taskID; // @[bbgemm.scala 203:44]
  wire [63:0] binaryOp_indvars_iv_next7934_io_Out_0_bits_data; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_Out_1_ready; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_Out_1_valid; // @[bbgemm.scala 203:44]
  wire [63:0] binaryOp_indvars_iv_next7934_io_Out_1_bits_data; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_LeftIO_ready; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_LeftIO_valid; // @[bbgemm.scala 203:44]
  wire [63:0] binaryOp_indvars_iv_next7934_io_LeftIO_bits_data; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_RightIO_ready; // @[bbgemm.scala 203:44]
  wire  binaryOp_indvars_iv_next7934_io_RightIO_valid; // @[bbgemm.scala 203:44]
  wire  icmp_exitcond8135_clock; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_reset; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_enable_ready; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_enable_valid; // @[bbgemm.scala 206:33]
  wire [4:0] icmp_exitcond8135_io_enable_bits_taskID; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_enable_bits_control; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_Out_0_ready; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_Out_0_valid; // @[bbgemm.scala 206:33]
  wire [4:0] icmp_exitcond8135_io_Out_0_bits_taskID; // @[bbgemm.scala 206:33]
  wire [63:0] icmp_exitcond8135_io_Out_0_bits_data; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_LeftIO_ready; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_LeftIO_valid; // @[bbgemm.scala 206:33]
  wire [63:0] icmp_exitcond8135_io_LeftIO_bits_data; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_RightIO_ready; // @[bbgemm.scala 206:33]
  wire  icmp_exitcond8135_io_RightIO_valid; // @[bbgemm.scala 206:33]
  wire  br_36_clock; // @[bbgemm.scala 209:21]
  wire  br_36_reset; // @[bbgemm.scala 209:21]
  wire  br_36_io_enable_ready; // @[bbgemm.scala 209:21]
  wire  br_36_io_enable_valid; // @[bbgemm.scala 209:21]
  wire [4:0] br_36_io_enable_bits_taskID; // @[bbgemm.scala 209:21]
  wire  br_36_io_enable_bits_control; // @[bbgemm.scala 209:21]
  wire  br_36_io_CmpIO_ready; // @[bbgemm.scala 209:21]
  wire  br_36_io_CmpIO_valid; // @[bbgemm.scala 209:21]
  wire [4:0] br_36_io_CmpIO_bits_taskID; // @[bbgemm.scala 209:21]
  wire [63:0] br_36_io_CmpIO_bits_data; // @[bbgemm.scala 209:21]
  wire  br_36_io_TrueOutput_0_ready; // @[bbgemm.scala 209:21]
  wire  br_36_io_TrueOutput_0_valid; // @[bbgemm.scala 209:21]
  wire  br_36_io_TrueOutput_0_bits_control; // @[bbgemm.scala 209:21]
  wire  br_36_io_FalseOutput_0_ready; // @[bbgemm.scala 209:21]
  wire  br_36_io_FalseOutput_0_valid; // @[bbgemm.scala 209:21]
  wire [4:0] br_36_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 209:21]
  wire  br_36_io_FalseOutput_0_bits_control; // @[bbgemm.scala 209:21]
  wire  binaryOp_indvars_iv_next8337_clock; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_reset; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_enable_ready; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_enable_valid; // @[bbgemm.scala 212:44]
  wire [4:0] binaryOp_indvars_iv_next8337_io_enable_bits_taskID; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_enable_bits_control; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_Out_0_ready; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_Out_0_valid; // @[bbgemm.scala 212:44]
  wire [4:0] binaryOp_indvars_iv_next8337_io_Out_0_bits_taskID; // @[bbgemm.scala 212:44]
  wire [63:0] binaryOp_indvars_iv_next8337_io_Out_0_bits_data; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_Out_1_ready; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_Out_1_valid; // @[bbgemm.scala 212:44]
  wire [63:0] binaryOp_indvars_iv_next8337_io_Out_1_bits_data; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_LeftIO_ready; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_LeftIO_valid; // @[bbgemm.scala 212:44]
  wire [63:0] binaryOp_indvars_iv_next8337_io_LeftIO_bits_data; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_RightIO_ready; // @[bbgemm.scala 212:44]
  wire  binaryOp_indvars_iv_next8337_io_RightIO_valid; // @[bbgemm.scala 212:44]
  wire  icmp_cmp238_clock; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_reset; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_enable_ready; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_enable_valid; // @[bbgemm.scala 215:27]
  wire [4:0] icmp_cmp238_io_enable_bits_taskID; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_enable_bits_control; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_Out_0_ready; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_Out_0_valid; // @[bbgemm.scala 215:27]
  wire [4:0] icmp_cmp238_io_Out_0_bits_taskID; // @[bbgemm.scala 215:27]
  wire [63:0] icmp_cmp238_io_Out_0_bits_data; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_LeftIO_ready; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_LeftIO_valid; // @[bbgemm.scala 215:27]
  wire [63:0] icmp_cmp238_io_LeftIO_bits_data; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_RightIO_ready; // @[bbgemm.scala 215:27]
  wire  icmp_cmp238_io_RightIO_valid; // @[bbgemm.scala 215:27]
  wire  br_39_clock; // @[bbgemm.scala 218:21]
  wire  br_39_reset; // @[bbgemm.scala 218:21]
  wire  br_39_io_enable_ready; // @[bbgemm.scala 218:21]
  wire  br_39_io_enable_valid; // @[bbgemm.scala 218:21]
  wire [4:0] br_39_io_enable_bits_taskID; // @[bbgemm.scala 218:21]
  wire  br_39_io_enable_bits_control; // @[bbgemm.scala 218:21]
  wire  br_39_io_CmpIO_ready; // @[bbgemm.scala 218:21]
  wire  br_39_io_CmpIO_valid; // @[bbgemm.scala 218:21]
  wire [4:0] br_39_io_CmpIO_bits_taskID; // @[bbgemm.scala 218:21]
  wire [63:0] br_39_io_CmpIO_bits_data; // @[bbgemm.scala 218:21]
  wire  br_39_io_TrueOutput_0_ready; // @[bbgemm.scala 218:21]
  wire  br_39_io_TrueOutput_0_valid; // @[bbgemm.scala 218:21]
  wire [4:0] br_39_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 218:21]
  wire  br_39_io_TrueOutput_0_bits_control; // @[bbgemm.scala 218:21]
  wire  br_39_io_FalseOutput_0_ready; // @[bbgemm.scala 218:21]
  wire  br_39_io_FalseOutput_0_valid; // @[bbgemm.scala 218:21]
  wire  br_39_io_FalseOutput_0_bits_control; // @[bbgemm.scala 218:21]
  wire  binaryOp_indvars_iv_next8540_clock; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_reset; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_enable_ready; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_enable_valid; // @[bbgemm.scala 221:44]
  wire [4:0] binaryOp_indvars_iv_next8540_io_enable_bits_taskID; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_enable_bits_control; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_Out_0_ready; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_Out_0_valid; // @[bbgemm.scala 221:44]
  wire [4:0] binaryOp_indvars_iv_next8540_io_Out_0_bits_taskID; // @[bbgemm.scala 221:44]
  wire [63:0] binaryOp_indvars_iv_next8540_io_Out_0_bits_data; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_Out_1_ready; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_Out_1_valid; // @[bbgemm.scala 221:44]
  wire [63:0] binaryOp_indvars_iv_next8540_io_Out_1_bits_data; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_LeftIO_ready; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_LeftIO_valid; // @[bbgemm.scala 221:44]
  wire [63:0] binaryOp_indvars_iv_next8540_io_LeftIO_bits_data; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_RightIO_ready; // @[bbgemm.scala 221:44]
  wire  binaryOp_indvars_iv_next8540_io_RightIO_valid; // @[bbgemm.scala 221:44]
  wire  icmp_cmp41_clock; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_reset; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_enable_ready; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_enable_valid; // @[bbgemm.scala 224:26]
  wire [4:0] icmp_cmp41_io_enable_bits_taskID; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_enable_bits_control; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_Out_0_ready; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_Out_0_valid; // @[bbgemm.scala 224:26]
  wire [4:0] icmp_cmp41_io_Out_0_bits_taskID; // @[bbgemm.scala 224:26]
  wire [63:0] icmp_cmp41_io_Out_0_bits_data; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_LeftIO_ready; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_LeftIO_valid; // @[bbgemm.scala 224:26]
  wire [63:0] icmp_cmp41_io_LeftIO_bits_data; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_RightIO_ready; // @[bbgemm.scala 224:26]
  wire  icmp_cmp41_io_RightIO_valid; // @[bbgemm.scala 224:26]
  wire  br_42_clock; // @[bbgemm.scala 227:21]
  wire  br_42_reset; // @[bbgemm.scala 227:21]
  wire  br_42_io_enable_ready; // @[bbgemm.scala 227:21]
  wire  br_42_io_enable_valid; // @[bbgemm.scala 227:21]
  wire [4:0] br_42_io_enable_bits_taskID; // @[bbgemm.scala 227:21]
  wire  br_42_io_enable_bits_control; // @[bbgemm.scala 227:21]
  wire  br_42_io_CmpIO_ready; // @[bbgemm.scala 227:21]
  wire  br_42_io_CmpIO_valid; // @[bbgemm.scala 227:21]
  wire [4:0] br_42_io_CmpIO_bits_taskID; // @[bbgemm.scala 227:21]
  wire [63:0] br_42_io_CmpIO_bits_data; // @[bbgemm.scala 227:21]
  wire  br_42_io_TrueOutput_0_ready; // @[bbgemm.scala 227:21]
  wire  br_42_io_TrueOutput_0_valid; // @[bbgemm.scala 227:21]
  wire [4:0] br_42_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 227:21]
  wire  br_42_io_TrueOutput_0_bits_control; // @[bbgemm.scala 227:21]
  wire  br_42_io_FalseOutput_0_ready; // @[bbgemm.scala 227:21]
  wire  br_42_io_FalseOutput_0_valid; // @[bbgemm.scala 227:21]
  wire  br_42_io_FalseOutput_0_bits_control; // @[bbgemm.scala 227:21]
  wire  ret_43_clock; // @[bbgemm.scala 230:22]
  wire  ret_43_reset; // @[bbgemm.scala 230:22]
  wire  ret_43_io_In_enable_ready; // @[bbgemm.scala 230:22]
  wire  ret_43_io_In_enable_valid; // @[bbgemm.scala 230:22]
  wire [4:0] ret_43_io_In_enable_bits_taskID; // @[bbgemm.scala 230:22]
  wire  ret_43_io_Out_ready; // @[bbgemm.scala 230:22]
  wire  ret_43_io_Out_valid; // @[bbgemm.scala 230:22]
  wire  const0_clock; // @[bbgemm.scala 239:22]
  wire  const0_reset; // @[bbgemm.scala 239:22]
  wire  const0_io_enable_ready; // @[bbgemm.scala 239:22]
  wire  const0_io_enable_valid; // @[bbgemm.scala 239:22]
  wire [4:0] const0_io_enable_bits_taskID; // @[bbgemm.scala 239:22]
  wire  const0_io_enable_bits_control; // @[bbgemm.scala 239:22]
  wire  const0_io_Out_ready; // @[bbgemm.scala 239:22]
  wire  const0_io_Out_valid; // @[bbgemm.scala 239:22]
  wire [4:0] const0_io_Out_bits_taskID; // @[bbgemm.scala 239:22]
  wire  const1_clock; // @[bbgemm.scala 242:22]
  wire  const1_reset; // @[bbgemm.scala 242:22]
  wire  const1_io_enable_ready; // @[bbgemm.scala 242:22]
  wire  const1_io_enable_valid; // @[bbgemm.scala 242:22]
  wire [4:0] const1_io_enable_bits_taskID; // @[bbgemm.scala 242:22]
  wire  const1_io_enable_bits_control; // @[bbgemm.scala 242:22]
  wire  const1_io_Out_ready; // @[bbgemm.scala 242:22]
  wire  const1_io_Out_valid; // @[bbgemm.scala 242:22]
  wire [4:0] const1_io_Out_bits_taskID; // @[bbgemm.scala 242:22]
  wire  const2_clock; // @[bbgemm.scala 245:22]
  wire  const2_reset; // @[bbgemm.scala 245:22]
  wire  const2_io_enable_ready; // @[bbgemm.scala 245:22]
  wire  const2_io_enable_valid; // @[bbgemm.scala 245:22]
  wire [4:0] const2_io_enable_bits_taskID; // @[bbgemm.scala 245:22]
  wire  const2_io_enable_bits_control; // @[bbgemm.scala 245:22]
  wire  const2_io_Out_ready; // @[bbgemm.scala 245:22]
  wire  const2_io_Out_valid; // @[bbgemm.scala 245:22]
  wire [4:0] const2_io_Out_bits_taskID; // @[bbgemm.scala 245:22]
  wire  const3_clock; // @[bbgemm.scala 248:22]
  wire  const3_reset; // @[bbgemm.scala 248:22]
  wire  const3_io_enable_ready; // @[bbgemm.scala 248:22]
  wire  const3_io_enable_valid; // @[bbgemm.scala 248:22]
  wire [4:0] const3_io_enable_bits_taskID; // @[bbgemm.scala 248:22]
  wire  const3_io_enable_bits_control; // @[bbgemm.scala 248:22]
  wire  const3_io_Out_ready; // @[bbgemm.scala 248:22]
  wire  const3_io_Out_valid; // @[bbgemm.scala 248:22]
  wire  const4_clock; // @[bbgemm.scala 251:22]
  wire  const4_reset; // @[bbgemm.scala 251:22]
  wire  const4_io_enable_ready; // @[bbgemm.scala 251:22]
  wire  const4_io_enable_valid; // @[bbgemm.scala 251:22]
  wire [4:0] const4_io_enable_bits_taskID; // @[bbgemm.scala 251:22]
  wire  const4_io_enable_bits_control; // @[bbgemm.scala 251:22]
  wire  const4_io_Out_ready; // @[bbgemm.scala 251:22]
  wire  const4_io_Out_valid; // @[bbgemm.scala 251:22]
  wire [4:0] const4_io_Out_bits_taskID; // @[bbgemm.scala 251:22]
  wire  const5_clock; // @[bbgemm.scala 254:22]
  wire  const5_reset; // @[bbgemm.scala 254:22]
  wire  const5_io_enable_ready; // @[bbgemm.scala 254:22]
  wire  const5_io_enable_valid; // @[bbgemm.scala 254:22]
  wire [4:0] const5_io_enable_bits_taskID; // @[bbgemm.scala 254:22]
  wire  const5_io_enable_bits_control; // @[bbgemm.scala 254:22]
  wire  const5_io_Out_ready; // @[bbgemm.scala 254:22]
  wire  const5_io_Out_valid; // @[bbgemm.scala 254:22]
  wire  const6_clock; // @[bbgemm.scala 257:22]
  wire  const6_reset; // @[bbgemm.scala 257:22]
  wire  const6_io_enable_ready; // @[bbgemm.scala 257:22]
  wire  const6_io_enable_valid; // @[bbgemm.scala 257:22]
  wire [4:0] const6_io_enable_bits_taskID; // @[bbgemm.scala 257:22]
  wire  const6_io_enable_bits_control; // @[bbgemm.scala 257:22]
  wire  const6_io_Out_ready; // @[bbgemm.scala 257:22]
  wire  const6_io_Out_valid; // @[bbgemm.scala 257:22]
  wire [4:0] const6_io_Out_bits_taskID; // @[bbgemm.scala 257:22]
  wire  const7_clock; // @[bbgemm.scala 260:22]
  wire  const7_reset; // @[bbgemm.scala 260:22]
  wire  const7_io_enable_ready; // @[bbgemm.scala 260:22]
  wire  const7_io_enable_valid; // @[bbgemm.scala 260:22]
  wire [4:0] const7_io_enable_bits_taskID; // @[bbgemm.scala 260:22]
  wire  const7_io_enable_bits_control; // @[bbgemm.scala 260:22]
  wire  const7_io_Out_ready; // @[bbgemm.scala 260:22]
  wire  const7_io_Out_valid; // @[bbgemm.scala 260:22]
  wire  const8_clock; // @[bbgemm.scala 263:22]
  wire  const8_reset; // @[bbgemm.scala 263:22]
  wire  const8_io_enable_ready; // @[bbgemm.scala 263:22]
  wire  const8_io_enable_valid; // @[bbgemm.scala 263:22]
  wire [4:0] const8_io_enable_bits_taskID; // @[bbgemm.scala 263:22]
  wire  const8_io_enable_bits_control; // @[bbgemm.scala 263:22]
  wire  const8_io_Out_ready; // @[bbgemm.scala 263:22]
  wire  const8_io_Out_valid; // @[bbgemm.scala 263:22]
  wire  const9_clock; // @[bbgemm.scala 266:22]
  wire  const9_reset; // @[bbgemm.scala 266:22]
  wire  const9_io_enable_ready; // @[bbgemm.scala 266:22]
  wire  const9_io_enable_valid; // @[bbgemm.scala 266:22]
  wire [4:0] const9_io_enable_bits_taskID; // @[bbgemm.scala 266:22]
  wire  const9_io_enable_bits_control; // @[bbgemm.scala 266:22]
  wire  const9_io_Out_ready; // @[bbgemm.scala 266:22]
  wire  const9_io_Out_valid; // @[bbgemm.scala 266:22]
  wire  const10_clock; // @[bbgemm.scala 269:23]
  wire  const10_reset; // @[bbgemm.scala 269:23]
  wire  const10_io_enable_ready; // @[bbgemm.scala 269:23]
  wire  const10_io_enable_valid; // @[bbgemm.scala 269:23]
  wire [4:0] const10_io_enable_bits_taskID; // @[bbgemm.scala 269:23]
  wire  const10_io_enable_bits_control; // @[bbgemm.scala 269:23]
  wire  const10_io_Out_ready; // @[bbgemm.scala 269:23]
  wire  const10_io_Out_valid; // @[bbgemm.scala 269:23]
  wire  const11_clock; // @[bbgemm.scala 272:23]
  wire  const11_reset; // @[bbgemm.scala 272:23]
  wire  const11_io_enable_ready; // @[bbgemm.scala 272:23]
  wire  const11_io_enable_valid; // @[bbgemm.scala 272:23]
  wire [4:0] const11_io_enable_bits_taskID; // @[bbgemm.scala 272:23]
  wire  const11_io_enable_bits_control; // @[bbgemm.scala 272:23]
  wire  const11_io_Out_ready; // @[bbgemm.scala 272:23]
  wire  const11_io_Out_valid; // @[bbgemm.scala 272:23]
  wire  const12_clock; // @[bbgemm.scala 275:23]
  wire  const12_reset; // @[bbgemm.scala 275:23]
  wire  const12_io_enable_ready; // @[bbgemm.scala 275:23]
  wire  const12_io_enable_valid; // @[bbgemm.scala 275:23]
  wire [4:0] const12_io_enable_bits_taskID; // @[bbgemm.scala 275:23]
  wire  const12_io_enable_bits_control; // @[bbgemm.scala 275:23]
  wire  const12_io_Out_ready; // @[bbgemm.scala 275:23]
  wire  const12_io_Out_valid; // @[bbgemm.scala 275:23]
  wire  const13_clock; // @[bbgemm.scala 278:23]
  wire  const13_reset; // @[bbgemm.scala 278:23]
  wire  const13_io_enable_ready; // @[bbgemm.scala 278:23]
  wire  const13_io_enable_valid; // @[bbgemm.scala 278:23]
  wire [4:0] const13_io_enable_bits_taskID; // @[bbgemm.scala 278:23]
  wire  const13_io_enable_bits_control; // @[bbgemm.scala 278:23]
  wire  const13_io_Out_ready; // @[bbgemm.scala 278:23]
  wire  const13_io_Out_valid; // @[bbgemm.scala 278:23]
  wire  const14_clock; // @[bbgemm.scala 281:23]
  wire  const14_reset; // @[bbgemm.scala 281:23]
  wire  const14_io_enable_ready; // @[bbgemm.scala 281:23]
  wire  const14_io_enable_valid; // @[bbgemm.scala 281:23]
  wire [4:0] const14_io_enable_bits_taskID; // @[bbgemm.scala 281:23]
  wire  const14_io_enable_bits_control; // @[bbgemm.scala 281:23]
  wire  const14_io_Out_ready; // @[bbgemm.scala 281:23]
  wire  const14_io_Out_valid; // @[bbgemm.scala 281:23]
  wire  const15_clock; // @[bbgemm.scala 284:23]
  wire  const15_reset; // @[bbgemm.scala 284:23]
  wire  const15_io_enable_ready; // @[bbgemm.scala 284:23]
  wire  const15_io_enable_valid; // @[bbgemm.scala 284:23]
  wire [4:0] const15_io_enable_bits_taskID; // @[bbgemm.scala 284:23]
  wire  const15_io_enable_bits_control; // @[bbgemm.scala 284:23]
  wire  const15_io_Out_ready; // @[bbgemm.scala 284:23]
  wire  const15_io_Out_valid; // @[bbgemm.scala 284:23]
  wire  const16_clock; // @[bbgemm.scala 287:23]
  wire  const16_reset; // @[bbgemm.scala 287:23]
  wire  const16_io_enable_ready; // @[bbgemm.scala 287:23]
  wire  const16_io_enable_valid; // @[bbgemm.scala 287:23]
  wire [4:0] const16_io_enable_bits_taskID; // @[bbgemm.scala 287:23]
  wire  const16_io_enable_bits_control; // @[bbgemm.scala 287:23]
  wire  const16_io_Out_ready; // @[bbgemm.scala 287:23]
  wire  const16_io_Out_valid; // @[bbgemm.scala 287:23]
  CacheMemoryEngine MemCtrl ( // @[bbgemm.scala 34:23]
    .clock(MemCtrl_clock),
    .reset(MemCtrl_reset),
    .io_rd_mem_0_MemReq_ready(MemCtrl_io_rd_mem_0_MemReq_ready),
    .io_rd_mem_0_MemReq_valid(MemCtrl_io_rd_mem_0_MemReq_valid),
    .io_rd_mem_0_MemReq_bits_addr(MemCtrl_io_rd_mem_0_MemReq_bits_addr),
    .io_rd_mem_0_MemResp_valid(MemCtrl_io_rd_mem_0_MemResp_valid),
    .io_rd_mem_0_MemResp_bits_data(MemCtrl_io_rd_mem_0_MemResp_bits_data),
    .io_rd_mem_1_MemReq_ready(MemCtrl_io_rd_mem_1_MemReq_ready),
    .io_rd_mem_1_MemReq_valid(MemCtrl_io_rd_mem_1_MemReq_valid),
    .io_rd_mem_1_MemReq_bits_addr(MemCtrl_io_rd_mem_1_MemReq_bits_addr),
    .io_rd_mem_1_MemResp_valid(MemCtrl_io_rd_mem_1_MemResp_valid),
    .io_rd_mem_1_MemResp_bits_data(MemCtrl_io_rd_mem_1_MemResp_bits_data),
    .io_rd_mem_2_MemReq_ready(MemCtrl_io_rd_mem_2_MemReq_ready),
    .io_rd_mem_2_MemReq_valid(MemCtrl_io_rd_mem_2_MemReq_valid),
    .io_rd_mem_2_MemReq_bits_addr(MemCtrl_io_rd_mem_2_MemReq_bits_addr),
    .io_rd_mem_2_MemResp_valid(MemCtrl_io_rd_mem_2_MemResp_valid),
    .io_rd_mem_2_MemResp_bits_data(MemCtrl_io_rd_mem_2_MemResp_bits_data),
    .io_wr_mem_0_MemReq_ready(MemCtrl_io_wr_mem_0_MemReq_ready),
    .io_wr_mem_0_MemReq_valid(MemCtrl_io_wr_mem_0_MemReq_valid),
    .io_wr_mem_0_MemReq_bits_addr(MemCtrl_io_wr_mem_0_MemReq_bits_addr),
    .io_wr_mem_0_MemReq_bits_data(MemCtrl_io_wr_mem_0_MemReq_bits_data),
    .io_wr_mem_0_MemResp_valid(MemCtrl_io_wr_mem_0_MemResp_valid),
    .io_cache_MemReq_ready(MemCtrl_io_cache_MemReq_ready),
    .io_cache_MemReq_valid(MemCtrl_io_cache_MemReq_valid),
    .io_cache_MemReq_bits_addr(MemCtrl_io_cache_MemReq_bits_addr),
    .io_cache_MemReq_bits_data(MemCtrl_io_cache_MemReq_bits_data),
    .io_cache_MemReq_bits_mask(MemCtrl_io_cache_MemReq_bits_mask),
    .io_cache_MemReq_bits_tag(MemCtrl_io_cache_MemReq_bits_tag),
    .io_cache_MemResp_valid(MemCtrl_io_cache_MemResp_valid),
    .io_cache_MemResp_bits_data(MemCtrl_io_cache_MemResp_bits_data),
    .io_cache_MemResp_bits_tag(MemCtrl_io_cache_MemResp_bits_tag)
  );
  SplitCallDCR ArgSplitter ( // @[bbgemm.scala 38:27]
    .clock(ArgSplitter_clock),
    .reset(ArgSplitter_reset),
    .io_In_ready(ArgSplitter_io_In_ready),
    .io_In_valid(ArgSplitter_io_In_valid),
    .io_In_bits_dataPtrs_field2_data(ArgSplitter_io_In_bits_dataPtrs_field2_data),
    .io_In_bits_dataPtrs_field1_data(ArgSplitter_io_In_bits_dataPtrs_field1_data),
    .io_In_bits_dataPtrs_field0_data(ArgSplitter_io_In_bits_dataPtrs_field0_data),
    .io_Out_enable_ready(ArgSplitter_io_Out_enable_ready),
    .io_Out_enable_valid(ArgSplitter_io_Out_enable_valid),
    .io_Out_enable_bits_control(ArgSplitter_io_Out_enable_bits_control),
    .io_Out_dataPtrs_field2_0_ready(ArgSplitter_io_Out_dataPtrs_field2_0_ready),
    .io_Out_dataPtrs_field2_0_valid(ArgSplitter_io_Out_dataPtrs_field2_0_valid),
    .io_Out_dataPtrs_field2_0_bits_data(ArgSplitter_io_Out_dataPtrs_field2_0_bits_data),
    .io_Out_dataPtrs_field1_0_ready(ArgSplitter_io_Out_dataPtrs_field1_0_ready),
    .io_Out_dataPtrs_field1_0_valid(ArgSplitter_io_Out_dataPtrs_field1_0_valid),
    .io_Out_dataPtrs_field1_0_bits_data(ArgSplitter_io_Out_dataPtrs_field1_0_bits_data),
    .io_Out_dataPtrs_field0_0_ready(ArgSplitter_io_Out_dataPtrs_field0_0_ready),
    .io_Out_dataPtrs_field0_0_valid(ArgSplitter_io_Out_dataPtrs_field0_0_valid),
    .io_Out_dataPtrs_field0_0_bits_data(ArgSplitter_io_Out_dataPtrs_field0_0_bits_data)
  );
  LoopBlockNode Loop_0 ( // @[bbgemm.scala 47:22]
    .clock(Loop_0_clock),
    .reset(Loop_0_reset),
    .io_enable_ready(Loop_0_io_enable_ready),
    .io_enable_valid(Loop_0_io_enable_valid),
    .io_enable_bits_taskID(Loop_0_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_0_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_0_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_0_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_0_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_0_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_0_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_0_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_0_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_0_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_0_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_0_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_0_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_0_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_0_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_0_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_data(Loop_0_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_0_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_0_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_0_io_InLiveIn_5_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_0_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_0_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_0_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field5_1_ready(Loop_0_io_OutLiveIn_field5_1_ready),
    .io_OutLiveIn_field5_1_valid(Loop_0_io_OutLiveIn_field5_1_valid),
    .io_OutLiveIn_field5_1_bits_data(Loop_0_io_OutLiveIn_field5_1_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_0_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_0_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_data(Loop_0_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_0_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_0_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_0_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_0_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_0_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_0_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_0_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_0_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_0_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_0_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_0_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_0_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_0_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_0_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_0_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_0_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_0_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_0_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_0_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_0_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_0_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_0_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_0_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_0_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_0_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_0_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_0_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_0_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_0_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_0_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_0_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_0_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_0_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_0_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_0_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_0_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_0_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_0_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_0_io_loopExit_0_bits_control)
  );
  LoopBlockNode_1 Loop_1 ( // @[bbgemm.scala 49:22]
    .clock(Loop_1_clock),
    .reset(Loop_1_reset),
    .io_enable_ready(Loop_1_io_enable_ready),
    .io_enable_valid(Loop_1_io_enable_valid),
    .io_enable_bits_taskID(Loop_1_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_1_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_1_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_1_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_1_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_1_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_1_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_1_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_1_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_1_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_1_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_1_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_1_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_1_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_1_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_1_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_data(Loop_1_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_1_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_1_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_1_io_InLiveIn_5_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_1_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_1_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_1_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_1_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_1_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_data(Loop_1_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field4_1_ready(Loop_1_io_OutLiveIn_field4_1_ready),
    .io_OutLiveIn_field4_1_valid(Loop_1_io_OutLiveIn_field4_1_valid),
    .io_OutLiveIn_field4_1_bits_data(Loop_1_io_OutLiveIn_field4_1_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_1_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_1_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_1_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_1_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_1_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_1_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_1_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_1_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_1_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_1_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_1_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_1_io_OutLiveIn_field0_0_bits_data),
    .io_OutLiveIn_field0_1_ready(Loop_1_io_OutLiveIn_field0_1_ready),
    .io_OutLiveIn_field0_1_valid(Loop_1_io_OutLiveIn_field0_1_valid),
    .io_OutLiveIn_field0_1_bits_data(Loop_1_io_OutLiveIn_field0_1_bits_data),
    .io_activate_loop_start_ready(Loop_1_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_1_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_1_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_1_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_1_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_1_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_1_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_1_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_1_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_1_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_1_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_1_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_1_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_1_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_1_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_1_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_1_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_1_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_1_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_1_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_1_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_1_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_1_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_1_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_1_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_1_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_1_io_loopExit_0_bits_control)
  );
  LoopBlockNode_2 Loop_2 ( // @[bbgemm.scala 51:22]
    .clock(Loop_2_clock),
    .reset(Loop_2_reset),
    .io_enable_ready(Loop_2_io_enable_ready),
    .io_enable_valid(Loop_2_io_enable_valid),
    .io_enable_bits_taskID(Loop_2_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_2_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_2_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_2_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_2_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_2_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_2_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_2_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_2_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_2_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_2_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_2_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_2_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_2_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_2_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_2_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_data(Loop_2_io_InLiveIn_4_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_2_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_2_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_data(Loop_2_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_2_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_2_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_2_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_2_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_2_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_2_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_2_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_2_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_2_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_2_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_2_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_2_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_2_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_2_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_2_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_2_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_2_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_2_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_2_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_2_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_2_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_2_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_2_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_2_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_2_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_2_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_2_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_2_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_2_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_2_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_2_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_2_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_2_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_2_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_2_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_2_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_2_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_2_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_2_io_loopExit_0_bits_control)
  );
  LoopBlockNode_3 Loop_3 ( // @[bbgemm.scala 53:22]
    .clock(Loop_3_clock),
    .reset(Loop_3_reset),
    .io_enable_ready(Loop_3_io_enable_ready),
    .io_enable_valid(Loop_3_io_enable_valid),
    .io_enable_bits_taskID(Loop_3_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_3_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_3_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_3_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_3_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_3_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_3_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_3_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_3_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_3_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_3_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_3_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_3_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_3_io_InLiveIn_3_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_3_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_3_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_3_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_3_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_3_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_3_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_3_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_3_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_3_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_3_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_3_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_3_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_3_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_3_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_3_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_3_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_3_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_3_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_3_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_3_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_3_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_3_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_3_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_3_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_3_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_3_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_3_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_3_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_3_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_3_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_3_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_3_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_3_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_3_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_3_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_3_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_3_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_3_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_3_io_loopExit_0_bits_control)
  );
  LoopBlockNode_4 Loop_4 ( // @[bbgemm.scala 55:22]
    .clock(Loop_4_clock),
    .reset(Loop_4_reset),
    .io_enable_ready(Loop_4_io_enable_ready),
    .io_enable_valid(Loop_4_io_enable_valid),
    .io_enable_bits_control(Loop_4_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_4_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_4_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_4_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_4_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_4_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_4_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_4_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_4_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_4_io_InLiveIn_2_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_4_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_4_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_4_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_4_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_4_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_4_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_4_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_4_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_4_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_4_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_4_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_4_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_4_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_4_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_4_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_4_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_4_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_4_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_4_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_4_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_4_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_4_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_4_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_4_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_4_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_4_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_4_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_4_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_4_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_4_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_4_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_4_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_4_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_4_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_4_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_4_io_loopExit_0_bits_control)
  );
  BasicBlockNoMaskFastNode bb_entry0 ( // @[bbgemm.scala 63:25]
    .clock(bb_entry0_clock),
    .reset(bb_entry0_reset),
    .io_predicateIn_0_ready(bb_entry0_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_entry0_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_control(bb_entry0_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_entry0_io_Out_0_ready),
    .io_Out_0_valid(bb_entry0_io_Out_0_valid),
    .io_Out_0_bits_control(bb_entry0_io_Out_0_bits_control)
  );
  BasicBlockNode bb_loopkk1 ( // @[bbgemm.scala 65:26]
    .clock(bb_loopkk1_clock),
    .reset(bb_loopkk1_reset),
    .io_MaskBB_0_ready(bb_loopkk1_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_loopkk1_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_loopkk1_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_loopkk1_io_Out_0_ready),
    .io_Out_0_valid(bb_loopkk1_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_loopkk1_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_loopkk1_io_Out_0_bits_control),
    .io_Out_1_ready(bb_loopkk1_io_Out_1_ready),
    .io_Out_1_valid(bb_loopkk1_io_Out_1_valid),
    .io_Out_1_bits_control(bb_loopkk1_io_Out_1_bits_control),
    .io_Out_2_ready(bb_loopkk1_io_Out_2_ready),
    .io_Out_2_valid(bb_loopkk1_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_loopkk1_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_loopkk1_io_Out_2_bits_control),
    .io_predicateIn_0_ready(bb_loopkk1_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_loopkk1_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_loopkk1_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_loopkk1_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_loopkk1_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_loopkk1_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_loopkk1_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_loopkk1_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_1 bb_loopi2 ( // @[bbgemm.scala 67:25]
    .clock(bb_loopi2_clock),
    .reset(bb_loopi2_reset),
    .io_MaskBB_0_ready(bb_loopi2_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_loopi2_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_loopi2_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_loopi2_io_Out_0_ready),
    .io_Out_0_valid(bb_loopi2_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_loopi2_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_loopi2_io_Out_0_bits_control),
    .io_Out_1_ready(bb_loopi2_io_Out_1_ready),
    .io_Out_1_valid(bb_loopi2_io_Out_1_valid),
    .io_Out_1_bits_control(bb_loopi2_io_Out_1_bits_control),
    .io_Out_2_ready(bb_loopi2_io_Out_2_ready),
    .io_Out_2_valid(bb_loopi2_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_loopi2_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_loopi2_io_Out_2_bits_control),
    .io_predicateIn_0_ready(bb_loopi2_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_loopi2_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_loopi2_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_loopi2_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_loopi2_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_loopi2_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_loopi2_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_loopi2_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_2 bb_loopk3 ( // @[bbgemm.scala 69:25]
    .clock(bb_loopk3_clock),
    .reset(bb_loopk3_reset),
    .io_MaskBB_0_ready(bb_loopk3_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_loopk3_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_loopk3_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_loopk3_io_Out_0_ready),
    .io_Out_0_valid(bb_loopk3_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_loopk3_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_loopk3_io_Out_0_bits_control),
    .io_Out_1_ready(bb_loopk3_io_Out_1_ready),
    .io_Out_1_valid(bb_loopk3_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_loopk3_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_loopk3_io_Out_1_bits_control),
    .io_Out_2_ready(bb_loopk3_io_Out_2_ready),
    .io_Out_2_valid(bb_loopk3_io_Out_2_valid),
    .io_Out_2_bits_control(bb_loopk3_io_Out_2_bits_control),
    .io_Out_3_ready(bb_loopk3_io_Out_3_ready),
    .io_Out_3_valid(bb_loopk3_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_loopk3_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_loopk3_io_Out_3_bits_control),
    .io_Out_4_ready(bb_loopk3_io_Out_4_ready),
    .io_Out_4_valid(bb_loopk3_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_loopk3_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_loopk3_io_Out_4_bits_control),
    .io_predicateIn_0_ready(bb_loopk3_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_loopk3_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_loopk3_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_loopk3_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_loopk3_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_loopk3_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_loopk3_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_loopk3_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_3 bb_for_body94 ( // @[bbgemm.scala 71:29]
    .clock(bb_for_body94_clock),
    .reset(bb_for_body94_reset),
    .io_MaskBB_0_ready(bb_for_body94_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body94_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body94_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body94_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body94_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body94_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_body94_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body94_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body94_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body94_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body94_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body94_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body94_io_Out_2_valid),
    .io_Out_2_bits_control(bb_for_body94_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body94_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body94_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body94_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_body94_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body94_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body94_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body94_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_body94_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_body94_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body94_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_body94_io_Out_5_bits_taskID),
    .io_Out_5_bits_control(bb_for_body94_io_Out_5_bits_control),
    .io_Out_6_ready(bb_for_body94_io_Out_6_ready),
    .io_Out_6_valid(bb_for_body94_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_body94_io_Out_6_bits_taskID),
    .io_Out_6_bits_control(bb_for_body94_io_Out_6_bits_control),
    .io_Out_7_ready(bb_for_body94_io_Out_7_ready),
    .io_Out_7_valid(bb_for_body94_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_body94_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_for_body94_io_Out_7_bits_control),
    .io_Out_8_ready(bb_for_body94_io_Out_8_ready),
    .io_Out_8_valid(bb_for_body94_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_for_body94_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_for_body94_io_Out_8_bits_control),
    .io_Out_9_ready(bb_for_body94_io_Out_9_ready),
    .io_Out_9_valid(bb_for_body94_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_for_body94_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_for_body94_io_Out_9_bits_control),
    .io_predicateIn_0_ready(bb_for_body94_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body94_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body94_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body94_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body94_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body94_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body94_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body94_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_4 bb_for_body165 ( // @[bbgemm.scala 73:30]
    .clock(bb_for_body165_clock),
    .reset(bb_for_body165_reset),
    .io_MaskBB_0_ready(bb_for_body165_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body165_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body165_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body165_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body165_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body165_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_body165_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body165_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body165_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body165_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body165_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body165_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body165_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body165_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body165_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body165_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body165_io_Out_3_valid),
    .io_Out_3_bits_control(bb_for_body165_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body165_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body165_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body165_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_body165_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_body165_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body165_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_body165_io_Out_5_bits_taskID),
    .io_Out_5_bits_control(bb_for_body165_io_Out_5_bits_control),
    .io_Out_6_ready(bb_for_body165_io_Out_6_ready),
    .io_Out_6_valid(bb_for_body165_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_body165_io_Out_6_bits_taskID),
    .io_Out_6_bits_control(bb_for_body165_io_Out_6_bits_control),
    .io_Out_7_ready(bb_for_body165_io_Out_7_ready),
    .io_Out_7_valid(bb_for_body165_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_body165_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_for_body165_io_Out_7_bits_control),
    .io_Out_8_ready(bb_for_body165_io_Out_8_ready),
    .io_Out_8_valid(bb_for_body165_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_for_body165_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_for_body165_io_Out_8_bits_control),
    .io_Out_9_ready(bb_for_body165_io_Out_9_ready),
    .io_Out_9_valid(bb_for_body165_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_for_body165_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_for_body165_io_Out_9_bits_control),
    .io_Out_10_ready(bb_for_body165_io_Out_10_ready),
    .io_Out_10_valid(bb_for_body165_io_Out_10_valid),
    .io_Out_10_bits_taskID(bb_for_body165_io_Out_10_bits_taskID),
    .io_Out_10_bits_control(bb_for_body165_io_Out_10_bits_control),
    .io_Out_11_ready(bb_for_body165_io_Out_11_ready),
    .io_Out_11_valid(bb_for_body165_io_Out_11_valid),
    .io_Out_11_bits_taskID(bb_for_body165_io_Out_11_bits_taskID),
    .io_Out_11_bits_control(bb_for_body165_io_Out_11_bits_control),
    .io_Out_12_ready(bb_for_body165_io_Out_12_ready),
    .io_Out_12_valid(bb_for_body165_io_Out_12_valid),
    .io_Out_12_bits_taskID(bb_for_body165_io_Out_12_bits_taskID),
    .io_Out_12_bits_control(bb_for_body165_io_Out_12_bits_control),
    .io_Out_13_ready(bb_for_body165_io_Out_13_ready),
    .io_Out_13_valid(bb_for_body165_io_Out_13_valid),
    .io_Out_13_bits_taskID(bb_for_body165_io_Out_13_bits_taskID),
    .io_Out_13_bits_control(bb_for_body165_io_Out_13_bits_control),
    .io_Out_14_ready(bb_for_body165_io_Out_14_ready),
    .io_Out_14_valid(bb_for_body165_io_Out_14_valid),
    .io_Out_14_bits_taskID(bb_for_body165_io_Out_14_bits_taskID),
    .io_Out_14_bits_control(bb_for_body165_io_Out_14_bits_control),
    .io_Out_15_ready(bb_for_body165_io_Out_15_ready),
    .io_Out_15_valid(bb_for_body165_io_Out_15_valid),
    .io_Out_15_bits_taskID(bb_for_body165_io_Out_15_bits_taskID),
    .io_Out_15_bits_control(bb_for_body165_io_Out_15_bits_control),
    .io_Out_16_ready(bb_for_body165_io_Out_16_ready),
    .io_Out_16_valid(bb_for_body165_io_Out_16_valid),
    .io_Out_16_bits_taskID(bb_for_body165_io_Out_16_bits_taskID),
    .io_Out_16_bits_control(bb_for_body165_io_Out_16_bits_control),
    .io_Out_17_ready(bb_for_body165_io_Out_17_ready),
    .io_Out_17_valid(bb_for_body165_io_Out_17_valid),
    .io_Out_17_bits_taskID(bb_for_body165_io_Out_17_bits_taskID),
    .io_Out_17_bits_control(bb_for_body165_io_Out_17_bits_control),
    .io_predicateIn_0_ready(bb_for_body165_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body165_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body165_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body165_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body165_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body165_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body165_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body165_io_predicateIn_1_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_for_inc276 ( // @[bbgemm.scala 75:29]
    .clock(bb_for_inc276_clock),
    .reset(bb_for_inc276_reset),
    .io_predicateIn_0_ready(bb_for_inc276_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_inc276_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_inc276_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_inc276_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_inc276_io_Out_0_ready),
    .io_Out_0_valid(bb_for_inc276_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_inc276_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_inc276_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_inc276_io_Out_1_ready),
    .io_Out_1_valid(bb_for_inc276_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_inc276_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_inc276_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_inc276_io_Out_2_ready),
    .io_Out_2_valid(bb_for_inc276_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_inc276_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_inc276_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_inc276_io_Out_3_ready),
    .io_Out_3_valid(bb_for_inc276_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_inc276_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_inc276_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_inc276_io_Out_4_ready),
    .io_Out_4_valid(bb_for_inc276_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_inc276_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_inc276_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_2 bb_for_inc307 ( // @[bbgemm.scala 77:29]
    .clock(bb_for_inc307_clock),
    .reset(bb_for_inc307_reset),
    .io_predicateIn_0_ready(bb_for_inc307_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_inc307_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_inc307_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_inc307_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_inc307_io_Out_0_ready),
    .io_Out_0_valid(bb_for_inc307_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_inc307_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_inc307_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_inc307_io_Out_1_ready),
    .io_Out_1_valid(bb_for_inc307_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_inc307_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_inc307_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_inc307_io_Out_2_ready),
    .io_Out_2_valid(bb_for_inc307_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_inc307_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_inc307_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_inc307_io_Out_3_ready),
    .io_Out_3_valid(bb_for_inc307_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_inc307_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_inc307_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_inc307_io_Out_4_ready),
    .io_Out_4_valid(bb_for_inc307_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_inc307_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_inc307_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_3 bb_for_inc338 ( // @[bbgemm.scala 79:29]
    .clock(bb_for_inc338_clock),
    .reset(bb_for_inc338_reset),
    .io_predicateIn_0_ready(bb_for_inc338_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_inc338_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_inc338_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_inc338_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_inc338_io_Out_0_ready),
    .io_Out_0_valid(bb_for_inc338_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_inc338_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_inc338_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_inc338_io_Out_1_ready),
    .io_Out_1_valid(bb_for_inc338_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_inc338_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_inc338_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_inc338_io_Out_2_ready),
    .io_Out_2_valid(bb_for_inc338_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_inc338_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_inc338_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_inc338_io_Out_3_ready),
    .io_Out_3_valid(bb_for_inc338_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_inc338_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_inc338_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_inc338_io_Out_4_ready),
    .io_Out_4_valid(bb_for_inc338_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_inc338_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_inc338_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_4 bb_for_inc369 ( // @[bbgemm.scala 81:29]
    .clock(bb_for_inc369_clock),
    .reset(bb_for_inc369_reset),
    .io_predicateIn_0_ready(bb_for_inc369_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_inc369_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_inc369_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_inc369_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_inc369_io_Out_0_ready),
    .io_Out_0_valid(bb_for_inc369_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_inc369_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_inc369_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_inc369_io_Out_1_ready),
    .io_Out_1_valid(bb_for_inc369_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_inc369_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_inc369_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_inc369_io_Out_2_ready),
    .io_Out_2_valid(bb_for_inc369_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_inc369_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_inc369_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_inc369_io_Out_3_ready),
    .io_Out_3_valid(bb_for_inc369_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_inc369_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_inc369_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_inc369_io_Out_4_ready),
    .io_Out_4_valid(bb_for_inc369_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_inc369_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_inc369_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_5 bb_for_end3810 ( // @[bbgemm.scala 83:30]
    .clock(bb_for_end3810_clock),
    .reset(bb_for_end3810_reset),
    .io_predicateIn_0_ready(bb_for_end3810_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_end3810_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_end3810_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_end3810_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_end3810_io_Out_0_ready),
    .io_Out_0_valid(bb_for_end3810_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_end3810_io_Out_0_bits_taskID)
  );
  UBranchNode br_0 ( // @[bbgemm.scala 92:20]
    .clock(br_0_clock),
    .reset(br_0_reset),
    .io_enable_ready(br_0_io_enable_ready),
    .io_enable_valid(br_0_io_enable_valid),
    .io_enable_bits_control(br_0_io_enable_bits_control),
    .io_Out_0_ready(br_0_io_Out_0_ready),
    .io_Out_0_valid(br_0_io_Out_0_valid),
    .io_Out_0_bits_control(br_0_io_Out_0_bits_control)
  );
  PhiFastNode phiindvars_iv841 ( // @[bbgemm.scala 95:32]
    .clock(phiindvars_iv841_clock),
    .reset(phiindvars_iv841_reset),
    .io_enable_ready(phiindvars_iv841_io_enable_ready),
    .io_enable_valid(phiindvars_iv841_io_enable_valid),
    .io_enable_bits_control(phiindvars_iv841_io_enable_bits_control),
    .io_InData_0_ready(phiindvars_iv841_io_InData_0_ready),
    .io_InData_0_valid(phiindvars_iv841_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiindvars_iv841_io_InData_0_bits_taskID),
    .io_InData_1_ready(phiindvars_iv841_io_InData_1_ready),
    .io_InData_1_valid(phiindvars_iv841_io_InData_1_valid),
    .io_InData_1_bits_taskID(phiindvars_iv841_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phiindvars_iv841_io_InData_1_bits_data),
    .io_Mask_ready(phiindvars_iv841_io_Mask_ready),
    .io_Mask_valid(phiindvars_iv841_io_Mask_valid),
    .io_Mask_bits(phiindvars_iv841_io_Mask_bits),
    .io_Out_0_ready(phiindvars_iv841_io_Out_0_ready),
    .io_Out_0_valid(phiindvars_iv841_io_Out_0_valid),
    .io_Out_0_bits_data(phiindvars_iv841_io_Out_0_bits_data),
    .io_Out_1_ready(phiindvars_iv841_io_Out_1_ready),
    .io_Out_1_valid(phiindvars_iv841_io_Out_1_valid),
    .io_Out_1_bits_data(phiindvars_iv841_io_Out_1_bits_data)
  );
  UBranchNode_1 br_2 ( // @[bbgemm.scala 97:20]
    .clock(br_2_clock),
    .reset(br_2_reset),
    .io_enable_ready(br_2_io_enable_ready),
    .io_enable_valid(br_2_io_enable_valid),
    .io_enable_bits_taskID(br_2_io_enable_bits_taskID),
    .io_enable_bits_control(br_2_io_enable_bits_control),
    .io_Out_0_ready(br_2_io_Out_0_ready),
    .io_Out_0_valid(br_2_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_2_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_2_io_Out_0_bits_control)
  );
  PhiFastNode_1 phiindvars_iv823 ( // @[bbgemm.scala 100:32]
    .clock(phiindvars_iv823_clock),
    .reset(phiindvars_iv823_reset),
    .io_enable_ready(phiindvars_iv823_io_enable_ready),
    .io_enable_valid(phiindvars_iv823_io_enable_valid),
    .io_enable_bits_control(phiindvars_iv823_io_enable_bits_control),
    .io_InData_0_ready(phiindvars_iv823_io_InData_0_ready),
    .io_InData_0_valid(phiindvars_iv823_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiindvars_iv823_io_InData_0_bits_taskID),
    .io_InData_1_ready(phiindvars_iv823_io_InData_1_ready),
    .io_InData_1_valid(phiindvars_iv823_io_InData_1_valid),
    .io_InData_1_bits_taskID(phiindvars_iv823_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phiindvars_iv823_io_InData_1_bits_data),
    .io_Mask_ready(phiindvars_iv823_io_Mask_ready),
    .io_Mask_valid(phiindvars_iv823_io_Mask_valid),
    .io_Mask_bits(phiindvars_iv823_io_Mask_bits),
    .io_Out_0_ready(phiindvars_iv823_io_Out_0_ready),
    .io_Out_0_valid(phiindvars_iv823_io_Out_0_valid),
    .io_Out_0_bits_data(phiindvars_iv823_io_Out_0_bits_data),
    .io_Out_1_ready(phiindvars_iv823_io_Out_1_ready),
    .io_Out_1_valid(phiindvars_iv823_io_Out_1_valid),
    .io_Out_1_bits_data(phiindvars_iv823_io_Out_1_bits_data)
  );
  UBranchNode_2 br_4 ( // @[bbgemm.scala 104:20]
    .clock(br_4_clock),
    .reset(br_4_reset),
    .io_enable_ready(br_4_io_enable_ready),
    .io_enable_valid(br_4_io_enable_valid),
    .io_enable_bits_taskID(br_4_io_enable_bits_taskID),
    .io_enable_bits_control(br_4_io_enable_bits_control),
    .io_Out_0_ready(br_4_io_Out_0_ready),
    .io_Out_0_valid(br_4_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_4_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_4_io_Out_0_bits_control)
  );
  PhiFastNode_2 phiindvars_iv785 ( // @[bbgemm.scala 107:32]
    .clock(phiindvars_iv785_clock),
    .reset(phiindvars_iv785_reset),
    .io_enable_ready(phiindvars_iv785_io_enable_ready),
    .io_enable_valid(phiindvars_iv785_io_enable_valid),
    .io_enable_bits_control(phiindvars_iv785_io_enable_bits_control),
    .io_InData_0_ready(phiindvars_iv785_io_InData_0_ready),
    .io_InData_0_valid(phiindvars_iv785_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiindvars_iv785_io_InData_0_bits_taskID),
    .io_InData_1_ready(phiindvars_iv785_io_InData_1_ready),
    .io_InData_1_valid(phiindvars_iv785_io_InData_1_valid),
    .io_InData_1_bits_taskID(phiindvars_iv785_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phiindvars_iv785_io_InData_1_bits_data),
    .io_Mask_ready(phiindvars_iv785_io_Mask_ready),
    .io_Mask_valid(phiindvars_iv785_io_Mask_valid),
    .io_Mask_bits(phiindvars_iv785_io_Mask_bits),
    .io_Out_0_ready(phiindvars_iv785_io_Out_0_ready),
    .io_Out_0_valid(phiindvars_iv785_io_Out_0_valid),
    .io_Out_0_bits_data(phiindvars_iv785_io_Out_0_bits_data),
    .io_Out_1_ready(phiindvars_iv785_io_Out_1_ready),
    .io_Out_1_valid(phiindvars_iv785_io_Out_1_valid),
    .io_Out_1_bits_data(phiindvars_iv785_io_Out_1_bits_data)
  );
  ComputeNode binaryOp_6 ( // @[bbgemm.scala 119:26]
    .clock(binaryOp_6_clock),
    .reset(binaryOp_6_reset),
    .io_enable_ready(binaryOp_6_io_enable_ready),
    .io_enable_valid(binaryOp_6_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_6_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_6_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_6_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_6_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_6_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_6_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_6_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_6_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_6_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_6_io_RightIO_valid)
  );
  UBranchNode_3 br_7 ( // @[bbgemm.scala 122:20]
    .clock(br_7_clock),
    .reset(br_7_reset),
    .io_enable_ready(br_7_io_enable_ready),
    .io_enable_valid(br_7_io_enable_valid),
    .io_enable_bits_taskID(br_7_io_enable_bits_taskID),
    .io_enable_bits_control(br_7_io_enable_bits_control),
    .io_Out_0_ready(br_7_io_Out_0_ready),
    .io_Out_0_valid(br_7_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_7_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_7_io_Out_0_bits_control)
  );
  PhiFastNode_3 phiindvars_iv718 ( // @[bbgemm.scala 125:32]
    .clock(phiindvars_iv718_clock),
    .reset(phiindvars_iv718_reset),
    .io_enable_ready(phiindvars_iv718_io_enable_ready),
    .io_enable_valid(phiindvars_iv718_io_enable_valid),
    .io_enable_bits_control(phiindvars_iv718_io_enable_bits_control),
    .io_InData_0_ready(phiindvars_iv718_io_InData_0_ready),
    .io_InData_0_valid(phiindvars_iv718_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiindvars_iv718_io_InData_0_bits_taskID),
    .io_InData_1_ready(phiindvars_iv718_io_InData_1_ready),
    .io_InData_1_valid(phiindvars_iv718_io_InData_1_valid),
    .io_InData_1_bits_taskID(phiindvars_iv718_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phiindvars_iv718_io_InData_1_bits_data),
    .io_Mask_ready(phiindvars_iv718_io_Mask_ready),
    .io_Mask_valid(phiindvars_iv718_io_Mask_valid),
    .io_Mask_bits(phiindvars_iv718_io_Mask_bits),
    .io_Out_0_ready(phiindvars_iv718_io_Out_0_ready),
    .io_Out_0_valid(phiindvars_iv718_io_Out_0_valid),
    .io_Out_0_bits_data(phiindvars_iv718_io_Out_0_bits_data),
    .io_Out_1_ready(phiindvars_iv718_io_Out_1_ready),
    .io_Out_1_valid(phiindvars_iv718_io_Out_1_valid),
    .io_Out_1_bits_data(phiindvars_iv718_io_Out_1_bits_data),
    .io_Out_2_ready(phiindvars_iv718_io_Out_2_ready),
    .io_Out_2_valid(phiindvars_iv718_io_Out_2_valid),
    .io_Out_2_bits_data(phiindvars_iv718_io_Out_2_bits_data)
  );
  ComputeNode_1 binaryOp_9 ( // @[bbgemm.scala 128:26]
    .clock(binaryOp_9_clock),
    .reset(binaryOp_9_reset),
    .io_enable_ready(binaryOp_9_io_enable_ready),
    .io_enable_valid(binaryOp_9_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_9_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_9_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_9_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_9_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_9_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_9_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_9_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_9_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_9_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_9_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_9_io_RightIO_bits_data)
  );
  ComputeNode_2 binaryOp_10 ( // @[bbgemm.scala 131:27]
    .clock(binaryOp_10_clock),
    .reset(binaryOp_10_reset),
    .io_enable_ready(binaryOp_10_io_enable_ready),
    .io_enable_valid(binaryOp_10_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_10_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_10_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_10_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_10_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_10_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_10_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_10_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_10_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_10_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_10_io_RightIO_valid)
  );
  ComputeNode_3 binaryOp_11 ( // @[bbgemm.scala 134:27]
    .clock(binaryOp_11_clock),
    .reset(binaryOp_11_reset),
    .io_enable_ready(binaryOp_11_io_enable_ready),
    .io_enable_valid(binaryOp_11_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_11_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_11_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_11_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_11_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_11_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_11_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_11_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_11_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_11_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_11_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_11_io_RightIO_bits_data)
  );
  ComputeNode_4 binaryOp_12 ( // @[bbgemm.scala 137:27]
    .clock(binaryOp_12_clock),
    .reset(binaryOp_12_reset),
    .io_enable_ready(binaryOp_12_io_enable_ready),
    .io_enable_valid(binaryOp_12_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_12_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_12_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_12_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_12_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_12_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_12_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_12_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_12_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_12_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_12_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_12_io_RightIO_bits_data)
  );
  GepNode Gep_arrayidx13 ( // @[bbgemm.scala 140:30]
    .clock(Gep_arrayidx13_clock),
    .reset(Gep_arrayidx13_reset),
    .io_enable_ready(Gep_arrayidx13_io_enable_ready),
    .io_enable_valid(Gep_arrayidx13_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx13_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx13_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx13_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx13_io_Out_0_valid),
    .io_Out_0_bits_data(Gep_arrayidx13_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx13_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx13_io_baseAddress_valid),
    .io_baseAddress_bits_data(Gep_arrayidx13_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx13_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx13_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx13_io_idx_0_bits_data)
  );
  UnTypLoadCache ld_14 ( // @[bbgemm.scala 143:21]
    .clock(ld_14_clock),
    .reset(ld_14_reset),
    .io_enable_ready(ld_14_io_enable_ready),
    .io_enable_valid(ld_14_io_enable_valid),
    .io_enable_bits_taskID(ld_14_io_enable_bits_taskID),
    .io_enable_bits_control(ld_14_io_enable_bits_control),
    .io_Out_0_ready(ld_14_io_Out_0_ready),
    .io_Out_0_valid(ld_14_io_Out_0_valid),
    .io_Out_0_bits_data(ld_14_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_14_io_GepAddr_ready),
    .io_GepAddr_valid(ld_14_io_GepAddr_valid),
    .io_GepAddr_bits_data(ld_14_io_GepAddr_bits_data),
    .io_MemReq_ready(ld_14_io_MemReq_ready),
    .io_MemReq_valid(ld_14_io_MemReq_valid),
    .io_MemReq_bits_addr(ld_14_io_MemReq_bits_addr),
    .io_MemResp_valid(ld_14_io_MemResp_valid),
    .io_MemResp_bits_data(ld_14_io_MemResp_bits_data)
  );
  UBranchNode_4 br_15 ( // @[bbgemm.scala 146:21]
    .clock(br_15_clock),
    .reset(br_15_reset),
    .io_enable_ready(br_15_io_enable_ready),
    .io_enable_valid(br_15_io_enable_valid),
    .io_enable_bits_taskID(br_15_io_enable_bits_taskID),
    .io_enable_bits_control(br_15_io_enable_bits_control),
    .io_Out_0_ready(br_15_io_Out_0_ready),
    .io_Out_0_valid(br_15_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_15_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_15_io_Out_0_bits_control)
  );
  PhiFastNode_4 phiindvars_iv16 ( // @[bbgemm.scala 149:31]
    .clock(phiindvars_iv16_clock),
    .reset(phiindvars_iv16_reset),
    .io_enable_ready(phiindvars_iv16_io_enable_ready),
    .io_enable_valid(phiindvars_iv16_io_enable_valid),
    .io_enable_bits_control(phiindvars_iv16_io_enable_bits_control),
    .io_InData_0_ready(phiindvars_iv16_io_InData_0_ready),
    .io_InData_0_valid(phiindvars_iv16_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiindvars_iv16_io_InData_0_bits_taskID),
    .io_InData_1_ready(phiindvars_iv16_io_InData_1_ready),
    .io_InData_1_valid(phiindvars_iv16_io_InData_1_valid),
    .io_InData_1_bits_taskID(phiindvars_iv16_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phiindvars_iv16_io_InData_1_bits_data),
    .io_Mask_ready(phiindvars_iv16_io_Mask_ready),
    .io_Mask_valid(phiindvars_iv16_io_Mask_valid),
    .io_Mask_bits(phiindvars_iv16_io_Mask_bits),
    .io_Out_0_ready(phiindvars_iv16_io_Out_0_ready),
    .io_Out_0_valid(phiindvars_iv16_io_Out_0_valid),
    .io_Out_0_bits_data(phiindvars_iv16_io_Out_0_bits_data),
    .io_Out_1_ready(phiindvars_iv16_io_Out_1_ready),
    .io_Out_1_valid(phiindvars_iv16_io_Out_1_valid),
    .io_Out_1_bits_data(phiindvars_iv16_io_Out_1_bits_data),
    .io_Out_2_ready(phiindvars_iv16_io_Out_2_ready),
    .io_Out_2_valid(phiindvars_iv16_io_Out_2_valid),
    .io_Out_2_bits_data(phiindvars_iv16_io_Out_2_bits_data)
  );
  ComputeNode_5 binaryOp_17 ( // @[bbgemm.scala 152:27]
    .clock(binaryOp_17_clock),
    .reset(binaryOp_17_reset),
    .io_enable_ready(binaryOp_17_io_enable_ready),
    .io_enable_valid(binaryOp_17_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_17_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_17_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_17_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_17_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_17_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_17_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_17_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_17_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_17_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_17_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_17_io_RightIO_bits_data)
  );
  ComputeNode_6 binaryOp_18 ( // @[bbgemm.scala 155:27]
    .clock(binaryOp_18_clock),
    .reset(binaryOp_18_reset),
    .io_enable_ready(binaryOp_18_io_enable_ready),
    .io_enable_valid(binaryOp_18_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_18_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_18_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_18_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_18_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_18_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_18_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_18_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_18_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_18_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_18_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_18_io_RightIO_bits_data)
  );
  GepNode_1 Gep_arrayidx2019 ( // @[bbgemm.scala 158:32]
    .clock(Gep_arrayidx2019_clock),
    .reset(Gep_arrayidx2019_reset),
    .io_enable_ready(Gep_arrayidx2019_io_enable_ready),
    .io_enable_valid(Gep_arrayidx2019_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx2019_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx2019_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx2019_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx2019_io_Out_0_valid),
    .io_Out_0_bits_data(Gep_arrayidx2019_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx2019_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx2019_io_baseAddress_valid),
    .io_baseAddress_bits_data(Gep_arrayidx2019_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx2019_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx2019_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx2019_io_idx_0_bits_data)
  );
  UnTypLoadCache_1 ld_20 ( // @[bbgemm.scala 161:21]
    .clock(ld_20_clock),
    .reset(ld_20_reset),
    .io_enable_ready(ld_20_io_enable_ready),
    .io_enable_valid(ld_20_io_enable_valid),
    .io_enable_bits_taskID(ld_20_io_enable_bits_taskID),
    .io_enable_bits_control(ld_20_io_enable_bits_control),
    .io_Out_0_ready(ld_20_io_Out_0_ready),
    .io_Out_0_valid(ld_20_io_Out_0_valid),
    .io_Out_0_bits_data(ld_20_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_20_io_GepAddr_ready),
    .io_GepAddr_valid(ld_20_io_GepAddr_valid),
    .io_GepAddr_bits_data(ld_20_io_GepAddr_bits_data),
    .io_MemReq_ready(ld_20_io_MemReq_ready),
    .io_MemReq_valid(ld_20_io_MemReq_valid),
    .io_MemReq_bits_addr(ld_20_io_MemReq_bits_addr),
    .io_MemResp_valid(ld_20_io_MemResp_valid),
    .io_MemResp_bits_data(ld_20_io_MemResp_bits_data)
  );
  FPComputeNode FP_mul2121 ( // @[bbgemm.scala 164:26]
    .clock(FP_mul2121_clock),
    .reset(FP_mul2121_reset),
    .io_enable_ready(FP_mul2121_io_enable_ready),
    .io_enable_valid(FP_mul2121_io_enable_valid),
    .io_enable_bits_taskID(FP_mul2121_io_enable_bits_taskID),
    .io_enable_bits_control(FP_mul2121_io_enable_bits_control),
    .io_Out_0_ready(FP_mul2121_io_Out_0_ready),
    .io_Out_0_valid(FP_mul2121_io_Out_0_valid),
    .io_Out_0_bits_data(FP_mul2121_io_Out_0_bits_data),
    .io_LeftIO_ready(FP_mul2121_io_LeftIO_ready),
    .io_LeftIO_valid(FP_mul2121_io_LeftIO_valid),
    .io_LeftIO_bits_data(FP_mul2121_io_LeftIO_bits_data),
    .io_RightIO_ready(FP_mul2121_io_RightIO_ready),
    .io_RightIO_valid(FP_mul2121_io_RightIO_valid),
    .io_RightIO_bits_data(FP_mul2121_io_RightIO_bits_data)
  );
  ComputeNode_7 binaryOp_22 ( // @[bbgemm.scala 167:27]
    .clock(binaryOp_22_clock),
    .reset(binaryOp_22_reset),
    .io_enable_ready(binaryOp_22_io_enable_ready),
    .io_enable_valid(binaryOp_22_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_22_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_22_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_22_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_22_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_22_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_22_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_22_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_22_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_22_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_22_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_22_io_RightIO_bits_data)
  );
  ComputeNode_8 binaryOp_23 ( // @[bbgemm.scala 170:27]
    .clock(binaryOp_23_clock),
    .reset(binaryOp_23_reset),
    .io_enable_ready(binaryOp_23_io_enable_ready),
    .io_enable_valid(binaryOp_23_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_23_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_23_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_23_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_23_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_23_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_23_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_23_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_23_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_23_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_23_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_23_io_RightIO_bits_data)
  );
  GepNode_2 Gep_arrayidx2524 ( // @[bbgemm.scala 173:32]
    .clock(Gep_arrayidx2524_clock),
    .reset(Gep_arrayidx2524_reset),
    .io_enable_ready(Gep_arrayidx2524_io_enable_ready),
    .io_enable_valid(Gep_arrayidx2524_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx2524_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx2524_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx2524_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx2524_io_Out_0_valid),
    .io_Out_0_bits_data(Gep_arrayidx2524_io_Out_0_bits_data),
    .io_Out_1_ready(Gep_arrayidx2524_io_Out_1_ready),
    .io_Out_1_valid(Gep_arrayidx2524_io_Out_1_valid),
    .io_Out_1_bits_data(Gep_arrayidx2524_io_Out_1_bits_data),
    .io_baseAddress_ready(Gep_arrayidx2524_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx2524_io_baseAddress_valid),
    .io_baseAddress_bits_data(Gep_arrayidx2524_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx2524_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx2524_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx2524_io_idx_0_bits_data)
  );
  UnTypLoadCache_2 ld_25 ( // @[bbgemm.scala 176:21]
    .clock(ld_25_clock),
    .reset(ld_25_reset),
    .io_enable_ready(ld_25_io_enable_ready),
    .io_enable_valid(ld_25_io_enable_valid),
    .io_enable_bits_taskID(ld_25_io_enable_bits_taskID),
    .io_enable_bits_control(ld_25_io_enable_bits_control),
    .io_Out_0_ready(ld_25_io_Out_0_ready),
    .io_Out_0_valid(ld_25_io_Out_0_valid),
    .io_Out_0_bits_data(ld_25_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_25_io_GepAddr_ready),
    .io_GepAddr_valid(ld_25_io_GepAddr_valid),
    .io_GepAddr_bits_data(ld_25_io_GepAddr_bits_data),
    .io_MemReq_ready(ld_25_io_MemReq_ready),
    .io_MemReq_valid(ld_25_io_MemReq_valid),
    .io_MemReq_bits_addr(ld_25_io_MemReq_bits_addr),
    .io_MemResp_valid(ld_25_io_MemResp_valid),
    .io_MemResp_bits_data(ld_25_io_MemResp_bits_data)
  );
  FPComputeNode_1 FP_add2626 ( // @[bbgemm.scala 179:26]
    .clock(FP_add2626_clock),
    .reset(FP_add2626_reset),
    .io_enable_ready(FP_add2626_io_enable_ready),
    .io_enable_valid(FP_add2626_io_enable_valid),
    .io_enable_bits_taskID(FP_add2626_io_enable_bits_taskID),
    .io_enable_bits_control(FP_add2626_io_enable_bits_control),
    .io_Out_0_ready(FP_add2626_io_Out_0_ready),
    .io_Out_0_valid(FP_add2626_io_Out_0_valid),
    .io_Out_0_bits_data(FP_add2626_io_Out_0_bits_data),
    .io_LeftIO_ready(FP_add2626_io_LeftIO_ready),
    .io_LeftIO_valid(FP_add2626_io_LeftIO_valid),
    .io_LeftIO_bits_data(FP_add2626_io_LeftIO_bits_data),
    .io_RightIO_ready(FP_add2626_io_RightIO_ready),
    .io_RightIO_valid(FP_add2626_io_RightIO_valid),
    .io_RightIO_bits_data(FP_add2626_io_RightIO_bits_data)
  );
  UnTypStoreCache st_27 ( // @[bbgemm.scala 182:21]
    .clock(st_27_clock),
    .reset(st_27_reset),
    .io_enable_ready(st_27_io_enable_ready),
    .io_enable_valid(st_27_io_enable_valid),
    .io_enable_bits_taskID(st_27_io_enable_bits_taskID),
    .io_enable_bits_control(st_27_io_enable_bits_control),
    .io_SuccOp_0_ready(st_27_io_SuccOp_0_ready),
    .io_SuccOp_0_valid(st_27_io_SuccOp_0_valid),
    .io_GepAddr_ready(st_27_io_GepAddr_ready),
    .io_GepAddr_valid(st_27_io_GepAddr_valid),
    .io_GepAddr_bits_data(st_27_io_GepAddr_bits_data),
    .io_inData_ready(st_27_io_inData_ready),
    .io_inData_valid(st_27_io_inData_valid),
    .io_inData_bits_data(st_27_io_inData_bits_data),
    .io_MemReq_ready(st_27_io_MemReq_ready),
    .io_MemReq_valid(st_27_io_MemReq_valid),
    .io_MemReq_bits_addr(st_27_io_MemReq_bits_addr),
    .io_MemReq_bits_data(st_27_io_MemReq_bits_data),
    .io_MemResp_valid(st_27_io_MemResp_valid)
  );
  ComputeNode_9 binaryOp_indvars_iv_next28 ( // @[bbgemm.scala 185:42]
    .clock(binaryOp_indvars_iv_next28_clock),
    .reset(binaryOp_indvars_iv_next28_reset),
    .io_enable_ready(binaryOp_indvars_iv_next28_io_enable_ready),
    .io_enable_valid(binaryOp_indvars_iv_next28_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_indvars_iv_next28_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_indvars_iv_next28_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_indvars_iv_next28_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_indvars_iv_next28_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_indvars_iv_next28_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_indvars_iv_next28_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_indvars_iv_next28_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_indvars_iv_next28_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_indvars_iv_next28_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_indvars_iv_next28_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_indvars_iv_next28_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_indvars_iv_next28_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_indvars_iv_next28_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_indvars_iv_next28_io_RightIO_valid)
  );
  ComputeNode_10 icmp_exitcond29 ( // @[bbgemm.scala 188:31]
    .clock(icmp_exitcond29_clock),
    .reset(icmp_exitcond29_reset),
    .io_enable_ready(icmp_exitcond29_io_enable_ready),
    .io_enable_valid(icmp_exitcond29_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond29_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond29_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond29_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond29_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond29_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond29_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond29_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond29_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond29_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond29_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond29_io_RightIO_valid)
  );
  CBranchNodeVariable br_30 ( // @[bbgemm.scala 191:21]
    .clock(br_30_clock),
    .reset(br_30_reset),
    .io_enable_ready(br_30_io_enable_ready),
    .io_enable_valid(br_30_io_enable_valid),
    .io_enable_bits_taskID(br_30_io_enable_bits_taskID),
    .io_enable_bits_control(br_30_io_enable_bits_control),
    .io_CmpIO_ready(br_30_io_CmpIO_ready),
    .io_CmpIO_valid(br_30_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_30_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_30_io_CmpIO_bits_data),
    .io_PredOp_0_ready(br_30_io_PredOp_0_ready),
    .io_PredOp_0_valid(br_30_io_PredOp_0_valid),
    .io_TrueOutput_0_ready(br_30_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_30_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_30_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_30_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_30_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_30_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_30_io_FalseOutput_0_bits_control)
  );
  ComputeNode_11 binaryOp_indvars_iv_next7231 ( // @[bbgemm.scala 194:44]
    .clock(binaryOp_indvars_iv_next7231_clock),
    .reset(binaryOp_indvars_iv_next7231_reset),
    .io_enable_ready(binaryOp_indvars_iv_next7231_io_enable_ready),
    .io_enable_valid(binaryOp_indvars_iv_next7231_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_indvars_iv_next7231_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_indvars_iv_next7231_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_indvars_iv_next7231_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_indvars_iv_next7231_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_indvars_iv_next7231_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_indvars_iv_next7231_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_indvars_iv_next7231_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_indvars_iv_next7231_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_indvars_iv_next7231_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_indvars_iv_next7231_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_indvars_iv_next7231_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_indvars_iv_next7231_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_indvars_iv_next7231_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_indvars_iv_next7231_io_RightIO_valid)
  );
  ComputeNode_12 icmp_exitcond7732 ( // @[bbgemm.scala 197:33]
    .clock(icmp_exitcond7732_clock),
    .reset(icmp_exitcond7732_reset),
    .io_enable_ready(icmp_exitcond7732_io_enable_ready),
    .io_enable_valid(icmp_exitcond7732_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond7732_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond7732_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond7732_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond7732_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond7732_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond7732_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond7732_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond7732_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond7732_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond7732_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond7732_io_RightIO_valid)
  );
  CBranchNodeVariable_1 br_33 ( // @[bbgemm.scala 200:21]
    .clock(br_33_clock),
    .reset(br_33_reset),
    .io_enable_ready(br_33_io_enable_ready),
    .io_enable_valid(br_33_io_enable_valid),
    .io_enable_bits_taskID(br_33_io_enable_bits_taskID),
    .io_enable_bits_control(br_33_io_enable_bits_control),
    .io_CmpIO_ready(br_33_io_CmpIO_ready),
    .io_CmpIO_valid(br_33_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_33_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_33_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_33_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_33_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_33_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_33_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_33_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_33_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_33_io_FalseOutput_0_bits_control)
  );
  ComputeNode_13 binaryOp_indvars_iv_next7934 ( // @[bbgemm.scala 203:44]
    .clock(binaryOp_indvars_iv_next7934_clock),
    .reset(binaryOp_indvars_iv_next7934_reset),
    .io_enable_ready(binaryOp_indvars_iv_next7934_io_enable_ready),
    .io_enable_valid(binaryOp_indvars_iv_next7934_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_indvars_iv_next7934_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_indvars_iv_next7934_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_indvars_iv_next7934_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_indvars_iv_next7934_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_indvars_iv_next7934_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_indvars_iv_next7934_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_indvars_iv_next7934_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_indvars_iv_next7934_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_indvars_iv_next7934_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_indvars_iv_next7934_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_indvars_iv_next7934_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_indvars_iv_next7934_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_indvars_iv_next7934_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_indvars_iv_next7934_io_RightIO_valid)
  );
  ComputeNode_14 icmp_exitcond8135 ( // @[bbgemm.scala 206:33]
    .clock(icmp_exitcond8135_clock),
    .reset(icmp_exitcond8135_reset),
    .io_enable_ready(icmp_exitcond8135_io_enable_ready),
    .io_enable_valid(icmp_exitcond8135_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond8135_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond8135_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond8135_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond8135_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond8135_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond8135_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond8135_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond8135_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond8135_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond8135_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond8135_io_RightIO_valid)
  );
  CBranchNodeVariable_2 br_36 ( // @[bbgemm.scala 209:21]
    .clock(br_36_clock),
    .reset(br_36_reset),
    .io_enable_ready(br_36_io_enable_ready),
    .io_enable_valid(br_36_io_enable_valid),
    .io_enable_bits_taskID(br_36_io_enable_bits_taskID),
    .io_enable_bits_control(br_36_io_enable_bits_control),
    .io_CmpIO_ready(br_36_io_CmpIO_ready),
    .io_CmpIO_valid(br_36_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_36_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_36_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_36_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_36_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_36_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_36_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_36_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_36_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_36_io_FalseOutput_0_bits_control)
  );
  ComputeNode_15 binaryOp_indvars_iv_next8337 ( // @[bbgemm.scala 212:44]
    .clock(binaryOp_indvars_iv_next8337_clock),
    .reset(binaryOp_indvars_iv_next8337_reset),
    .io_enable_ready(binaryOp_indvars_iv_next8337_io_enable_ready),
    .io_enable_valid(binaryOp_indvars_iv_next8337_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_indvars_iv_next8337_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_indvars_iv_next8337_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_indvars_iv_next8337_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_indvars_iv_next8337_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_indvars_iv_next8337_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_indvars_iv_next8337_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_indvars_iv_next8337_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_indvars_iv_next8337_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_indvars_iv_next8337_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_indvars_iv_next8337_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_indvars_iv_next8337_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_indvars_iv_next8337_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_indvars_iv_next8337_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_indvars_iv_next8337_io_RightIO_valid)
  );
  ComputeNode_16 icmp_cmp238 ( // @[bbgemm.scala 215:27]
    .clock(icmp_cmp238_clock),
    .reset(icmp_cmp238_reset),
    .io_enable_ready(icmp_cmp238_io_enable_ready),
    .io_enable_valid(icmp_cmp238_io_enable_valid),
    .io_enable_bits_taskID(icmp_cmp238_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_cmp238_io_enable_bits_control),
    .io_Out_0_ready(icmp_cmp238_io_Out_0_ready),
    .io_Out_0_valid(icmp_cmp238_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_cmp238_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_cmp238_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_cmp238_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_cmp238_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_cmp238_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_cmp238_io_RightIO_ready),
    .io_RightIO_valid(icmp_cmp238_io_RightIO_valid)
  );
  CBranchNodeVariable_3 br_39 ( // @[bbgemm.scala 218:21]
    .clock(br_39_clock),
    .reset(br_39_reset),
    .io_enable_ready(br_39_io_enable_ready),
    .io_enable_valid(br_39_io_enable_valid),
    .io_enable_bits_taskID(br_39_io_enable_bits_taskID),
    .io_enable_bits_control(br_39_io_enable_bits_control),
    .io_CmpIO_ready(br_39_io_CmpIO_ready),
    .io_CmpIO_valid(br_39_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_39_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_39_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_39_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_39_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_39_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_39_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_39_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_39_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_control(br_39_io_FalseOutput_0_bits_control)
  );
  ComputeNode_17 binaryOp_indvars_iv_next8540 ( // @[bbgemm.scala 221:44]
    .clock(binaryOp_indvars_iv_next8540_clock),
    .reset(binaryOp_indvars_iv_next8540_reset),
    .io_enable_ready(binaryOp_indvars_iv_next8540_io_enable_ready),
    .io_enable_valid(binaryOp_indvars_iv_next8540_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_indvars_iv_next8540_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_indvars_iv_next8540_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_indvars_iv_next8540_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_indvars_iv_next8540_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_indvars_iv_next8540_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_indvars_iv_next8540_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_indvars_iv_next8540_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_indvars_iv_next8540_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_indvars_iv_next8540_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_indvars_iv_next8540_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_indvars_iv_next8540_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_indvars_iv_next8540_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_indvars_iv_next8540_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_indvars_iv_next8540_io_RightIO_valid)
  );
  ComputeNode_18 icmp_cmp41 ( // @[bbgemm.scala 224:26]
    .clock(icmp_cmp41_clock),
    .reset(icmp_cmp41_reset),
    .io_enable_ready(icmp_cmp41_io_enable_ready),
    .io_enable_valid(icmp_cmp41_io_enable_valid),
    .io_enable_bits_taskID(icmp_cmp41_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_cmp41_io_enable_bits_control),
    .io_Out_0_ready(icmp_cmp41_io_Out_0_ready),
    .io_Out_0_valid(icmp_cmp41_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_cmp41_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_cmp41_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_cmp41_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_cmp41_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_cmp41_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_cmp41_io_RightIO_ready),
    .io_RightIO_valid(icmp_cmp41_io_RightIO_valid)
  );
  CBranchNodeVariable_4 br_42 ( // @[bbgemm.scala 227:21]
    .clock(br_42_clock),
    .reset(br_42_reset),
    .io_enable_ready(br_42_io_enable_ready),
    .io_enable_valid(br_42_io_enable_valid),
    .io_enable_bits_taskID(br_42_io_enable_bits_taskID),
    .io_enable_bits_control(br_42_io_enable_bits_control),
    .io_CmpIO_ready(br_42_io_CmpIO_ready),
    .io_CmpIO_valid(br_42_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_42_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_42_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_42_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_42_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_42_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_42_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_42_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_42_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_control(br_42_io_FalseOutput_0_bits_control)
  );
  RetNode2 ret_43 ( // @[bbgemm.scala 230:22]
    .clock(ret_43_clock),
    .reset(ret_43_reset),
    .io_In_enable_ready(ret_43_io_In_enable_ready),
    .io_In_enable_valid(ret_43_io_In_enable_valid),
    .io_In_enable_bits_taskID(ret_43_io_In_enable_bits_taskID),
    .io_Out_ready(ret_43_io_Out_ready),
    .io_Out_valid(ret_43_io_Out_valid)
  );
  ConstFastNode const0 ( // @[bbgemm.scala 239:22]
    .clock(const0_clock),
    .reset(const0_reset),
    .io_enable_ready(const0_io_enable_ready),
    .io_enable_valid(const0_io_enable_valid),
    .io_enable_bits_taskID(const0_io_enable_bits_taskID),
    .io_enable_bits_control(const0_io_enable_bits_control),
    .io_Out_ready(const0_io_Out_ready),
    .io_Out_valid(const0_io_Out_valid),
    .io_Out_bits_taskID(const0_io_Out_bits_taskID)
  );
  ConstFastNode const1 ( // @[bbgemm.scala 242:22]
    .clock(const1_clock),
    .reset(const1_reset),
    .io_enable_ready(const1_io_enable_ready),
    .io_enable_valid(const1_io_enable_valid),
    .io_enable_bits_taskID(const1_io_enable_bits_taskID),
    .io_enable_bits_control(const1_io_enable_bits_control),
    .io_Out_ready(const1_io_Out_ready),
    .io_Out_valid(const1_io_Out_valid),
    .io_Out_bits_taskID(const1_io_Out_bits_taskID)
  );
  ConstFastNode const2 ( // @[bbgemm.scala 245:22]
    .clock(const2_clock),
    .reset(const2_reset),
    .io_enable_ready(const2_io_enable_ready),
    .io_enable_valid(const2_io_enable_valid),
    .io_enable_bits_taskID(const2_io_enable_bits_taskID),
    .io_enable_bits_control(const2_io_enable_bits_control),
    .io_Out_ready(const2_io_Out_ready),
    .io_Out_valid(const2_io_Out_valid),
    .io_Out_bits_taskID(const2_io_Out_bits_taskID)
  );
  ConstFastNode_3 const3 ( // @[bbgemm.scala 248:22]
    .clock(const3_clock),
    .reset(const3_reset),
    .io_enable_ready(const3_io_enable_ready),
    .io_enable_valid(const3_io_enable_valid),
    .io_enable_bits_taskID(const3_io_enable_bits_taskID),
    .io_enable_bits_control(const3_io_enable_bits_control),
    .io_Out_ready(const3_io_Out_ready),
    .io_Out_valid(const3_io_Out_valid)
  );
  ConstFastNode const4 ( // @[bbgemm.scala 251:22]
    .clock(const4_clock),
    .reset(const4_reset),
    .io_enable_ready(const4_io_enable_ready),
    .io_enable_valid(const4_io_enable_valid),
    .io_enable_bits_taskID(const4_io_enable_bits_taskID),
    .io_enable_bits_control(const4_io_enable_bits_control),
    .io_Out_ready(const4_io_Out_ready),
    .io_Out_valid(const4_io_Out_valid),
    .io_Out_bits_taskID(const4_io_Out_bits_taskID)
  );
  ConstFastNode_3 const5 ( // @[bbgemm.scala 254:22]
    .clock(const5_clock),
    .reset(const5_reset),
    .io_enable_ready(const5_io_enable_ready),
    .io_enable_valid(const5_io_enable_valid),
    .io_enable_bits_taskID(const5_io_enable_bits_taskID),
    .io_enable_bits_control(const5_io_enable_bits_control),
    .io_Out_ready(const5_io_Out_ready),
    .io_Out_valid(const5_io_Out_valid)
  );
  ConstFastNode const6 ( // @[bbgemm.scala 257:22]
    .clock(const6_clock),
    .reset(const6_reset),
    .io_enable_ready(const6_io_enable_ready),
    .io_enable_valid(const6_io_enable_valid),
    .io_enable_bits_taskID(const6_io_enable_bits_taskID),
    .io_enable_bits_control(const6_io_enable_bits_control),
    .io_Out_ready(const6_io_Out_ready),
    .io_Out_valid(const6_io_Out_valid),
    .io_Out_bits_taskID(const6_io_Out_bits_taskID)
  );
  ConstFastNode_7 const7 ( // @[bbgemm.scala 260:22]
    .clock(const7_clock),
    .reset(const7_reset),
    .io_enable_ready(const7_io_enable_ready),
    .io_enable_valid(const7_io_enable_valid),
    .io_enable_bits_taskID(const7_io_enable_bits_taskID),
    .io_enable_bits_control(const7_io_enable_bits_control),
    .io_Out_ready(const7_io_Out_ready),
    .io_Out_valid(const7_io_Out_valid)
  );
  ConstFastNode_8 const8 ( // @[bbgemm.scala 263:22]
    .clock(const8_clock),
    .reset(const8_reset),
    .io_enable_ready(const8_io_enable_ready),
    .io_enable_valid(const8_io_enable_valid),
    .io_enable_bits_taskID(const8_io_enable_bits_taskID),
    .io_enable_bits_control(const8_io_enable_bits_control),
    .io_Out_ready(const8_io_Out_ready),
    .io_Out_valid(const8_io_Out_valid)
  );
  ConstFastNode_7 const9 ( // @[bbgemm.scala 266:22]
    .clock(const9_clock),
    .reset(const9_reset),
    .io_enable_ready(const9_io_enable_ready),
    .io_enable_valid(const9_io_enable_valid),
    .io_enable_bits_taskID(const9_io_enable_bits_taskID),
    .io_enable_bits_control(const9_io_enable_bits_control),
    .io_Out_ready(const9_io_Out_ready),
    .io_Out_valid(const9_io_Out_valid)
  );
  ConstFastNode_8 const10 ( // @[bbgemm.scala 269:23]
    .clock(const10_clock),
    .reset(const10_reset),
    .io_enable_ready(const10_io_enable_ready),
    .io_enable_valid(const10_io_enable_valid),
    .io_enable_bits_taskID(const10_io_enable_bits_taskID),
    .io_enable_bits_control(const10_io_enable_bits_control),
    .io_Out_ready(const10_io_Out_ready),
    .io_Out_valid(const10_io_Out_valid)
  );
  ConstFastNode_7 const11 ( // @[bbgemm.scala 272:23]
    .clock(const11_clock),
    .reset(const11_reset),
    .io_enable_ready(const11_io_enable_ready),
    .io_enable_valid(const11_io_enable_valid),
    .io_enable_bits_taskID(const11_io_enable_bits_taskID),
    .io_enable_bits_control(const11_io_enable_bits_control),
    .io_Out_ready(const11_io_Out_ready),
    .io_Out_valid(const11_io_Out_valid)
  );
  ConstFastNode_12 const12 ( // @[bbgemm.scala 275:23]
    .clock(const12_clock),
    .reset(const12_reset),
    .io_enable_ready(const12_io_enable_ready),
    .io_enable_valid(const12_io_enable_valid),
    .io_enable_bits_taskID(const12_io_enable_bits_taskID),
    .io_enable_bits_control(const12_io_enable_bits_control),
    .io_Out_ready(const12_io_Out_ready),
    .io_Out_valid(const12_io_Out_valid)
  );
  ConstFastNode_8 const13 ( // @[bbgemm.scala 278:23]
    .clock(const13_clock),
    .reset(const13_reset),
    .io_enable_ready(const13_io_enable_ready),
    .io_enable_valid(const13_io_enable_valid),
    .io_enable_bits_taskID(const13_io_enable_bits_taskID),
    .io_enable_bits_control(const13_io_enable_bits_control),
    .io_Out_ready(const13_io_Out_ready),
    .io_Out_valid(const13_io_Out_valid)
  );
  ConstFastNode_12 const14 ( // @[bbgemm.scala 281:23]
    .clock(const14_clock),
    .reset(const14_reset),
    .io_enable_ready(const14_io_enable_ready),
    .io_enable_valid(const14_io_enable_valid),
    .io_enable_bits_taskID(const14_io_enable_bits_taskID),
    .io_enable_bits_control(const14_io_enable_bits_control),
    .io_Out_ready(const14_io_Out_ready),
    .io_Out_valid(const14_io_Out_valid)
  );
  ConstFastNode_8 const15 ( // @[bbgemm.scala 284:23]
    .clock(const15_clock),
    .reset(const15_reset),
    .io_enable_ready(const15_io_enable_ready),
    .io_enable_valid(const15_io_enable_valid),
    .io_enable_bits_taskID(const15_io_enable_bits_taskID),
    .io_enable_bits_control(const15_io_enable_bits_control),
    .io_Out_ready(const15_io_Out_ready),
    .io_Out_valid(const15_io_Out_valid)
  );
  ConstFastNode_12 const16 ( // @[bbgemm.scala 287:23]
    .clock(const16_clock),
    .reset(const16_reset),
    .io_enable_ready(const16_io_enable_ready),
    .io_enable_valid(const16_io_enable_valid),
    .io_enable_bits_taskID(const16_io_enable_bits_taskID),
    .io_enable_bits_control(const16_io_enable_bits_control),
    .io_Out_ready(const16_io_Out_ready),
    .io_Out_valid(const16_io_Out_valid)
  );
  assign io_in_ready = ArgSplitter_io_In_ready; // @[bbgemm.scala 39:21]
  assign io_MemReq_valid = MemCtrl_io_cache_MemReq_valid; // @[bbgemm.scala 36:13]
  assign io_MemReq_bits_addr = MemCtrl_io_cache_MemReq_bits_addr; // @[bbgemm.scala 36:13]
  assign io_MemReq_bits_data = MemCtrl_io_cache_MemReq_bits_data; // @[bbgemm.scala 36:13]
  assign io_MemReq_bits_mask = MemCtrl_io_cache_MemReq_bits_mask; // @[bbgemm.scala 36:13]
  assign io_MemReq_bits_tag = MemCtrl_io_cache_MemReq_bits_tag; // @[bbgemm.scala 36:13]
  assign io_out_valid = ret_43_io_Out_valid; // @[bbgemm.scala 854:10]
  assign MemCtrl_clock = clock;
  assign MemCtrl_reset = reset;
  assign MemCtrl_io_rd_mem_0_MemReq_valid = ld_14_io_MemReq_valid; // @[bbgemm.scala 707:31]
  assign MemCtrl_io_rd_mem_0_MemReq_bits_addr = ld_14_io_MemReq_bits_addr; // @[bbgemm.scala 707:31]
  assign MemCtrl_io_rd_mem_1_MemReq_valid = ld_20_io_MemReq_valid; // @[bbgemm.scala 711:31]
  assign MemCtrl_io_rd_mem_1_MemReq_bits_addr = ld_20_io_MemReq_bits_addr; // @[bbgemm.scala 711:31]
  assign MemCtrl_io_rd_mem_2_MemReq_valid = ld_25_io_MemReq_valid; // @[bbgemm.scala 715:31]
  assign MemCtrl_io_rd_mem_2_MemReq_bits_addr = ld_25_io_MemReq_bits_addr; // @[bbgemm.scala 715:31]
  assign MemCtrl_io_wr_mem_0_MemReq_valid = st_27_io_MemReq_valid; // @[bbgemm.scala 719:31]
  assign MemCtrl_io_wr_mem_0_MemReq_bits_addr = st_27_io_MemReq_bits_addr; // @[bbgemm.scala 719:31]
  assign MemCtrl_io_wr_mem_0_MemReq_bits_data = st_27_io_MemReq_bits_data; // @[bbgemm.scala 719:31]
  assign MemCtrl_io_cache_MemReq_ready = io_MemReq_ready; // @[bbgemm.scala 36:13]
  assign MemCtrl_io_cache_MemResp_valid = io_MemResp_valid; // @[bbgemm.scala 37:28]
  assign MemCtrl_io_cache_MemResp_bits_data = io_MemResp_bits_data; // @[bbgemm.scala 37:28]
  assign MemCtrl_io_cache_MemResp_bits_tag = io_MemResp_bits_tag; // @[bbgemm.scala 37:28]
  assign ArgSplitter_clock = clock;
  assign ArgSplitter_reset = reset;
  assign ArgSplitter_io_In_valid = io_in_valid; // @[bbgemm.scala 39:21]
  assign ArgSplitter_io_In_bits_dataPtrs_field2_data = {{32'd0}, io_in_bits_dataPtrs_field2_data}; // @[bbgemm.scala 39:21]
  assign ArgSplitter_io_In_bits_dataPtrs_field1_data = {{32'd0}, io_in_bits_dataPtrs_field1_data}; // @[bbgemm.scala 39:21]
  assign ArgSplitter_io_In_bits_dataPtrs_field0_data = {{32'd0}, io_in_bits_dataPtrs_field0_data}; // @[bbgemm.scala 39:21]
  assign ArgSplitter_io_Out_enable_ready = bb_entry0_io_predicateIn_0_ready; // @[bbgemm.scala 295:31]
  assign ArgSplitter_io_Out_dataPtrs_field2_0_ready = Loop_4_io_InLiveIn_2_ready; // @[bbgemm.scala 433:25]
  assign ArgSplitter_io_Out_dataPtrs_field1_0_ready = Loop_4_io_InLiveIn_1_ready; // @[bbgemm.scala 431:25]
  assign ArgSplitter_io_Out_dataPtrs_field0_0_ready = Loop_4_io_InLiveIn_0_ready; // @[bbgemm.scala 429:25]
  assign Loop_0_clock = clock;
  assign Loop_0_reset = reset;
  assign Loop_0_io_enable_valid = br_15_io_Out_0_valid; // @[bbgemm.scala 345:20]
  assign Loop_0_io_enable_bits_taskID = br_15_io_Out_0_bits_taskID; // @[bbgemm.scala 345:20]
  assign Loop_0_io_enable_bits_control = br_15_io_Out_0_bits_control; // @[bbgemm.scala 345:20]
  assign Loop_0_io_InLiveIn_0_valid = binaryOp_10_io_Out_0_valid; // @[bbgemm.scala 387:25]
  assign Loop_0_io_InLiveIn_0_bits_data = binaryOp_10_io_Out_0_bits_data; // @[bbgemm.scala 387:25]
  assign Loop_0_io_InLiveIn_1_valid = ld_14_io_Out_0_valid; // @[bbgemm.scala 389:25]
  assign Loop_0_io_InLiveIn_1_bits_data = ld_14_io_Out_0_bits_data; // @[bbgemm.scala 389:25]
  assign Loop_0_io_InLiveIn_2_valid = Loop_1_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 391:25]
  assign Loop_0_io_InLiveIn_2_bits_data = Loop_1_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 391:25]
  assign Loop_0_io_InLiveIn_3_valid = Loop_1_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 393:25]
  assign Loop_0_io_InLiveIn_3_bits_data = Loop_1_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 393:25]
  assign Loop_0_io_InLiveIn_4_valid = Loop_1_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 395:25]
  assign Loop_0_io_InLiveIn_4_bits_data = Loop_1_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 395:25]
  assign Loop_0_io_InLiveIn_5_valid = Loop_1_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 397:25]
  assign Loop_0_io_InLiveIn_5_bits_data = Loop_1_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 397:25]
  assign Loop_0_io_OutLiveIn_field5_0_ready = binaryOp_17_io_RightIO_ready; // @[bbgemm.scala 451:26]
  assign Loop_0_io_OutLiveIn_field5_1_ready = binaryOp_22_io_RightIO_ready; // @[bbgemm.scala 453:26]
  assign Loop_0_io_OutLiveIn_field4_0_ready = Gep_arrayidx2524_io_baseAddress_ready; // @[bbgemm.scala 449:35]
  assign Loop_0_io_OutLiveIn_field3_0_ready = binaryOp_23_io_RightIO_ready; // @[bbgemm.scala 447:26]
  assign Loop_0_io_OutLiveIn_field2_0_ready = Gep_arrayidx2019_io_baseAddress_ready; // @[bbgemm.scala 445:35]
  assign Loop_0_io_OutLiveIn_field1_0_ready = FP_mul2121_io_LeftIO_ready; // @[bbgemm.scala 443:24]
  assign Loop_0_io_OutLiveIn_field0_0_ready = binaryOp_18_io_RightIO_ready; // @[bbgemm.scala 441:26]
  assign Loop_0_io_activate_loop_start_ready = bb_for_body165_io_predicateIn_1_ready; // @[bbgemm.scala 319:36]
  assign Loop_0_io_activate_loop_back_ready = bb_for_body165_io_predicateIn_0_ready; // @[bbgemm.scala 321:36]
  assign Loop_0_io_loopBack_0_valid = br_30_io_FalseOutput_0_valid; // @[bbgemm.scala 347:25]
  assign Loop_0_io_loopBack_0_bits_taskID = br_30_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 347:25]
  assign Loop_0_io_loopBack_0_bits_control = br_30_io_FalseOutput_0_bits_control; // @[bbgemm.scala 347:25]
  assign Loop_0_io_loopFinish_0_valid = br_30_io_TrueOutput_0_valid; // @[bbgemm.scala 349:27]
  assign Loop_0_io_loopFinish_0_bits_control = br_30_io_TrueOutput_0_bits_control; // @[bbgemm.scala 349:27]
  assign Loop_0_io_CarryDepenIn_0_valid = binaryOp_indvars_iv_next28_io_Out_0_valid; // @[bbgemm.scala 481:29]
  assign Loop_0_io_CarryDepenIn_0_bits_taskID = binaryOp_indvars_iv_next28_io_Out_0_bits_taskID; // @[bbgemm.scala 481:29]
  assign Loop_0_io_CarryDepenIn_0_bits_data = binaryOp_indvars_iv_next28_io_Out_0_bits_data; // @[bbgemm.scala 481:29]
  assign Loop_0_io_CarryDepenOut_field0_0_ready = phiindvars_iv16_io_InData_1_ready; // @[bbgemm.scala 497:32]
  assign Loop_0_io_loopExit_0_ready = bb_for_inc276_io_predicateIn_0_ready; // @[bbgemm.scala 323:35]
  assign Loop_1_clock = clock;
  assign Loop_1_reset = reset;
  assign Loop_1_io_enable_valid = br_7_io_Out_0_valid; // @[bbgemm.scala 351:20]
  assign Loop_1_io_enable_bits_taskID = br_7_io_Out_0_bits_taskID; // @[bbgemm.scala 351:20]
  assign Loop_1_io_enable_bits_control = br_7_io_Out_0_bits_control; // @[bbgemm.scala 351:20]
  assign Loop_1_io_InLiveIn_0_valid = binaryOp_6_io_Out_0_valid; // @[bbgemm.scala 399:25]
  assign Loop_1_io_InLiveIn_0_bits_data = binaryOp_6_io_Out_0_bits_data; // @[bbgemm.scala 399:25]
  assign Loop_1_io_InLiveIn_1_valid = Loop_2_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 401:25]
  assign Loop_1_io_InLiveIn_1_bits_data = Loop_2_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 401:25]
  assign Loop_1_io_InLiveIn_2_valid = Loop_2_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 403:25]
  assign Loop_1_io_InLiveIn_2_bits_data = Loop_2_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 403:25]
  assign Loop_1_io_InLiveIn_3_valid = Loop_2_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 405:25]
  assign Loop_1_io_InLiveIn_3_bits_data = Loop_2_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 405:25]
  assign Loop_1_io_InLiveIn_4_valid = Loop_2_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 407:25]
  assign Loop_1_io_InLiveIn_4_bits_data = Loop_2_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 407:25]
  assign Loop_1_io_InLiveIn_5_valid = Loop_2_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 409:25]
  assign Loop_1_io_InLiveIn_5_bits_data = Loop_2_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 409:25]
  assign Loop_1_io_OutLiveIn_field5_0_ready = Gep_arrayidx13_io_baseAddress_ready; // @[bbgemm.scala 461:33]
  assign Loop_1_io_OutLiveIn_field4_0_ready = binaryOp_9_io_RightIO_ready; // @[bbgemm.scala 457:25]
  assign Loop_1_io_OutLiveIn_field4_1_ready = binaryOp_11_io_RightIO_ready; // @[bbgemm.scala 459:26]
  assign Loop_1_io_OutLiveIn_field3_0_ready = Loop_0_io_InLiveIn_5_ready; // @[bbgemm.scala 397:25]
  assign Loop_1_io_OutLiveIn_field2_0_ready = Loop_0_io_InLiveIn_4_ready; // @[bbgemm.scala 395:25]
  assign Loop_1_io_OutLiveIn_field1_0_ready = Loop_0_io_InLiveIn_2_ready; // @[bbgemm.scala 391:25]
  assign Loop_1_io_OutLiveIn_field0_0_ready = Loop_0_io_InLiveIn_3_ready; // @[bbgemm.scala 393:25]
  assign Loop_1_io_OutLiveIn_field0_1_ready = binaryOp_12_io_RightIO_ready; // @[bbgemm.scala 455:26]
  assign Loop_1_io_activate_loop_start_ready = bb_for_body94_io_predicateIn_1_ready; // @[bbgemm.scala 315:35]
  assign Loop_1_io_activate_loop_back_ready = bb_for_body94_io_predicateIn_0_ready; // @[bbgemm.scala 317:35]
  assign Loop_1_io_loopBack_0_valid = br_33_io_FalseOutput_0_valid; // @[bbgemm.scala 353:25]
  assign Loop_1_io_loopBack_0_bits_taskID = br_33_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 353:25]
  assign Loop_1_io_loopBack_0_bits_control = br_33_io_FalseOutput_0_bits_control; // @[bbgemm.scala 353:25]
  assign Loop_1_io_loopFinish_0_valid = br_33_io_TrueOutput_0_valid; // @[bbgemm.scala 355:27]
  assign Loop_1_io_loopFinish_0_bits_control = br_33_io_TrueOutput_0_bits_control; // @[bbgemm.scala 355:27]
  assign Loop_1_io_CarryDepenIn_0_valid = binaryOp_indvars_iv_next7231_io_Out_0_valid; // @[bbgemm.scala 483:29]
  assign Loop_1_io_CarryDepenIn_0_bits_taskID = binaryOp_indvars_iv_next7231_io_Out_0_bits_taskID; // @[bbgemm.scala 483:29]
  assign Loop_1_io_CarryDepenIn_0_bits_data = binaryOp_indvars_iv_next7231_io_Out_0_bits_data; // @[bbgemm.scala 483:29]
  assign Loop_1_io_CarryDepenOut_field0_0_ready = phiindvars_iv718_io_InData_1_ready; // @[bbgemm.scala 499:33]
  assign Loop_1_io_loopExit_0_ready = bb_for_inc307_io_predicateIn_0_ready; // @[bbgemm.scala 325:35]
  assign Loop_2_clock = clock;
  assign Loop_2_reset = reset;
  assign Loop_2_io_enable_valid = br_4_io_Out_0_valid; // @[bbgemm.scala 357:20]
  assign Loop_2_io_enable_bits_taskID = br_4_io_Out_0_bits_taskID; // @[bbgemm.scala 357:20]
  assign Loop_2_io_enable_bits_control = br_4_io_Out_0_bits_control; // @[bbgemm.scala 357:20]
  assign Loop_2_io_InLiveIn_0_valid = phiindvars_iv823_io_Out_0_valid; // @[bbgemm.scala 411:25]
  assign Loop_2_io_InLiveIn_0_bits_data = phiindvars_iv823_io_Out_0_bits_data; // @[bbgemm.scala 411:25]
  assign Loop_2_io_InLiveIn_1_valid = Loop_3_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 413:25]
  assign Loop_2_io_InLiveIn_1_bits_data = Loop_3_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 413:25]
  assign Loop_2_io_InLiveIn_2_valid = Loop_3_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 415:25]
  assign Loop_2_io_InLiveIn_2_bits_data = Loop_3_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 415:25]
  assign Loop_2_io_InLiveIn_3_valid = Loop_3_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 417:25]
  assign Loop_2_io_InLiveIn_3_bits_data = Loop_3_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 417:25]
  assign Loop_2_io_InLiveIn_4_valid = Loop_3_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 419:25]
  assign Loop_2_io_InLiveIn_4_bits_data = Loop_3_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 419:25]
  assign Loop_2_io_OutLiveIn_field4_0_ready = Loop_1_io_InLiveIn_3_ready; // @[bbgemm.scala 405:25]
  assign Loop_2_io_OutLiveIn_field3_0_ready = Loop_1_io_InLiveIn_2_ready; // @[bbgemm.scala 403:25]
  assign Loop_2_io_OutLiveIn_field2_0_ready = Loop_1_io_InLiveIn_5_ready; // @[bbgemm.scala 409:25]
  assign Loop_2_io_OutLiveIn_field1_0_ready = Loop_1_io_InLiveIn_1_ready; // @[bbgemm.scala 401:25]
  assign Loop_2_io_OutLiveIn_field0_0_ready = Loop_1_io_InLiveIn_4_ready; // @[bbgemm.scala 407:25]
  assign Loop_2_io_activate_loop_start_ready = bb_loopk3_io_predicateIn_1_ready; // @[bbgemm.scala 311:31]
  assign Loop_2_io_activate_loop_back_ready = bb_loopk3_io_predicateIn_0_ready; // @[bbgemm.scala 313:31]
  assign Loop_2_io_loopBack_0_valid = br_36_io_FalseOutput_0_valid; // @[bbgemm.scala 359:25]
  assign Loop_2_io_loopBack_0_bits_taskID = br_36_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 359:25]
  assign Loop_2_io_loopBack_0_bits_control = br_36_io_FalseOutput_0_bits_control; // @[bbgemm.scala 359:25]
  assign Loop_2_io_loopFinish_0_valid = br_36_io_TrueOutput_0_valid; // @[bbgemm.scala 361:27]
  assign Loop_2_io_loopFinish_0_bits_control = br_36_io_TrueOutput_0_bits_control; // @[bbgemm.scala 361:27]
  assign Loop_2_io_CarryDepenIn_0_valid = binaryOp_indvars_iv_next7934_io_Out_0_valid; // @[bbgemm.scala 485:29]
  assign Loop_2_io_CarryDepenIn_0_bits_taskID = binaryOp_indvars_iv_next7934_io_Out_0_bits_taskID; // @[bbgemm.scala 485:29]
  assign Loop_2_io_CarryDepenIn_0_bits_data = binaryOp_indvars_iv_next7934_io_Out_0_bits_data; // @[bbgemm.scala 485:29]
  assign Loop_2_io_CarryDepenOut_field0_0_ready = phiindvars_iv785_io_InData_1_ready; // @[bbgemm.scala 501:33]
  assign Loop_2_io_loopExit_0_ready = bb_for_inc338_io_predicateIn_0_ready; // @[bbgemm.scala 327:35]
  assign Loop_3_clock = clock;
  assign Loop_3_reset = reset;
  assign Loop_3_io_enable_valid = br_2_io_Out_0_valid; // @[bbgemm.scala 363:20]
  assign Loop_3_io_enable_bits_taskID = br_2_io_Out_0_bits_taskID; // @[bbgemm.scala 363:20]
  assign Loop_3_io_enable_bits_control = br_2_io_Out_0_bits_control; // @[bbgemm.scala 363:20]
  assign Loop_3_io_InLiveIn_0_valid = phiindvars_iv841_io_Out_0_valid; // @[bbgemm.scala 421:25]
  assign Loop_3_io_InLiveIn_0_bits_data = phiindvars_iv841_io_Out_0_bits_data; // @[bbgemm.scala 421:25]
  assign Loop_3_io_InLiveIn_1_valid = Loop_4_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 423:25]
  assign Loop_3_io_InLiveIn_1_bits_data = Loop_4_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 423:25]
  assign Loop_3_io_InLiveIn_2_valid = Loop_4_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 425:25]
  assign Loop_3_io_InLiveIn_2_bits_data = Loop_4_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 425:25]
  assign Loop_3_io_InLiveIn_3_valid = Loop_4_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 427:25]
  assign Loop_3_io_InLiveIn_3_bits_data = Loop_4_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 427:25]
  assign Loop_3_io_OutLiveIn_field3_0_ready = Loop_2_io_InLiveIn_3_ready; // @[bbgemm.scala 417:25]
  assign Loop_3_io_OutLiveIn_field2_0_ready = Loop_2_io_InLiveIn_2_ready; // @[bbgemm.scala 415:25]
  assign Loop_3_io_OutLiveIn_field1_0_ready = Loop_2_io_InLiveIn_1_ready; // @[bbgemm.scala 413:25]
  assign Loop_3_io_OutLiveIn_field0_0_ready = Loop_2_io_InLiveIn_4_ready; // @[bbgemm.scala 419:25]
  assign Loop_3_io_activate_loop_start_ready = bb_loopi2_io_predicateIn_0_ready; // @[bbgemm.scala 307:31]
  assign Loop_3_io_activate_loop_back_ready = bb_loopi2_io_predicateIn_1_ready; // @[bbgemm.scala 309:31]
  assign Loop_3_io_loopBack_0_valid = br_39_io_TrueOutput_0_valid; // @[bbgemm.scala 365:25]
  assign Loop_3_io_loopBack_0_bits_taskID = br_39_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 365:25]
  assign Loop_3_io_loopBack_0_bits_control = br_39_io_TrueOutput_0_bits_control; // @[bbgemm.scala 365:25]
  assign Loop_3_io_loopFinish_0_valid = br_39_io_FalseOutput_0_valid; // @[bbgemm.scala 367:27]
  assign Loop_3_io_loopFinish_0_bits_control = br_39_io_FalseOutput_0_bits_control; // @[bbgemm.scala 367:27]
  assign Loop_3_io_CarryDepenIn_0_valid = binaryOp_indvars_iv_next8337_io_Out_0_valid; // @[bbgemm.scala 487:29]
  assign Loop_3_io_CarryDepenIn_0_bits_taskID = binaryOp_indvars_iv_next8337_io_Out_0_bits_taskID; // @[bbgemm.scala 487:29]
  assign Loop_3_io_CarryDepenIn_0_bits_data = binaryOp_indvars_iv_next8337_io_Out_0_bits_data; // @[bbgemm.scala 487:29]
  assign Loop_3_io_CarryDepenOut_field0_0_ready = phiindvars_iv823_io_InData_1_ready; // @[bbgemm.scala 503:33]
  assign Loop_3_io_loopExit_0_ready = bb_for_inc369_io_predicateIn_0_ready; // @[bbgemm.scala 329:35]
  assign Loop_4_clock = clock;
  assign Loop_4_reset = reset;
  assign Loop_4_io_enable_valid = br_0_io_Out_0_valid; // @[bbgemm.scala 369:20]
  assign Loop_4_io_enable_bits_control = br_0_io_Out_0_bits_control; // @[bbgemm.scala 369:20]
  assign Loop_4_io_InLiveIn_0_valid = ArgSplitter_io_Out_dataPtrs_field0_0_valid; // @[bbgemm.scala 429:25]
  assign Loop_4_io_InLiveIn_0_bits_data = ArgSplitter_io_Out_dataPtrs_field0_0_bits_data; // @[bbgemm.scala 429:25]
  assign Loop_4_io_InLiveIn_1_valid = ArgSplitter_io_Out_dataPtrs_field1_0_valid; // @[bbgemm.scala 431:25]
  assign Loop_4_io_InLiveIn_1_bits_data = ArgSplitter_io_Out_dataPtrs_field1_0_bits_data; // @[bbgemm.scala 431:25]
  assign Loop_4_io_InLiveIn_2_valid = ArgSplitter_io_Out_dataPtrs_field2_0_valid; // @[bbgemm.scala 433:25]
  assign Loop_4_io_InLiveIn_2_bits_data = ArgSplitter_io_Out_dataPtrs_field2_0_bits_data; // @[bbgemm.scala 433:25]
  assign Loop_4_io_OutLiveIn_field2_0_ready = Loop_3_io_InLiveIn_3_ready; // @[bbgemm.scala 427:25]
  assign Loop_4_io_OutLiveIn_field1_0_ready = Loop_3_io_InLiveIn_1_ready; // @[bbgemm.scala 423:25]
  assign Loop_4_io_OutLiveIn_field0_0_ready = Loop_3_io_InLiveIn_2_ready; // @[bbgemm.scala 425:25]
  assign Loop_4_io_activate_loop_start_ready = bb_loopkk1_io_predicateIn_0_ready; // @[bbgemm.scala 303:32]
  assign Loop_4_io_activate_loop_back_ready = bb_loopkk1_io_predicateIn_1_ready; // @[bbgemm.scala 305:32]
  assign Loop_4_io_loopBack_0_valid = br_42_io_TrueOutput_0_valid; // @[bbgemm.scala 371:25]
  assign Loop_4_io_loopBack_0_bits_taskID = br_42_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 371:25]
  assign Loop_4_io_loopBack_0_bits_control = br_42_io_TrueOutput_0_bits_control; // @[bbgemm.scala 371:25]
  assign Loop_4_io_loopFinish_0_valid = br_42_io_FalseOutput_0_valid; // @[bbgemm.scala 373:27]
  assign Loop_4_io_loopFinish_0_bits_control = br_42_io_FalseOutput_0_bits_control; // @[bbgemm.scala 373:27]
  assign Loop_4_io_CarryDepenIn_0_valid = binaryOp_indvars_iv_next8540_io_Out_0_valid; // @[bbgemm.scala 489:29]
  assign Loop_4_io_CarryDepenIn_0_bits_taskID = binaryOp_indvars_iv_next8540_io_Out_0_bits_taskID; // @[bbgemm.scala 489:29]
  assign Loop_4_io_CarryDepenIn_0_bits_data = binaryOp_indvars_iv_next8540_io_Out_0_bits_data; // @[bbgemm.scala 489:29]
  assign Loop_4_io_CarryDepenOut_field0_0_ready = phiindvars_iv841_io_InData_1_ready; // @[bbgemm.scala 505:33]
  assign Loop_4_io_loopExit_0_ready = bb_for_end3810_io_predicateIn_0_ready; // @[bbgemm.scala 331:36]
  assign bb_entry0_clock = clock;
  assign bb_entry0_reset = reset;
  assign bb_entry0_io_predicateIn_0_valid = ArgSplitter_io_Out_enable_valid; // @[bbgemm.scala 295:31]
  assign bb_entry0_io_predicateIn_0_bits_control = ArgSplitter_io_Out_enable_bits_control; // @[bbgemm.scala 295:31]
  assign bb_entry0_io_Out_0_ready = br_0_io_enable_ready; // @[bbgemm.scala 513:18]
  assign bb_loopkk1_clock = clock;
  assign bb_loopkk1_reset = reset;
  assign bb_loopkk1_io_MaskBB_0_ready = phiindvars_iv841_io_Mask_ready; // @[bbgemm.scala 685:28]
  assign bb_loopkk1_io_Out_0_ready = const0_io_enable_ready; // @[bbgemm.scala 516:20]
  assign bb_loopkk1_io_Out_1_ready = phiindvars_iv841_io_enable_ready; // @[bbgemm.scala 518:30]
  assign bb_loopkk1_io_Out_2_ready = br_2_io_enable_ready; // @[bbgemm.scala 521:18]
  assign bb_loopkk1_io_predicateIn_0_valid = Loop_4_io_activate_loop_start_valid; // @[bbgemm.scala 303:32]
  assign bb_loopkk1_io_predicateIn_0_bits_taskID = Loop_4_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 303:32]
  assign bb_loopkk1_io_predicateIn_0_bits_control = Loop_4_io_activate_loop_start_bits_control; // @[bbgemm.scala 303:32]
  assign bb_loopkk1_io_predicateIn_1_valid = Loop_4_io_activate_loop_back_valid; // @[bbgemm.scala 305:32]
  assign bb_loopkk1_io_predicateIn_1_bits_taskID = Loop_4_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 305:32]
  assign bb_loopkk1_io_predicateIn_1_bits_control = Loop_4_io_activate_loop_back_bits_control; // @[bbgemm.scala 305:32]
  assign bb_loopi2_clock = clock;
  assign bb_loopi2_reset = reset;
  assign bb_loopi2_io_MaskBB_0_ready = phiindvars_iv823_io_Mask_ready; // @[bbgemm.scala 687:28]
  assign bb_loopi2_io_Out_0_ready = const1_io_enable_ready; // @[bbgemm.scala 524:20]
  assign bb_loopi2_io_Out_1_ready = phiindvars_iv823_io_enable_ready; // @[bbgemm.scala 526:30]
  assign bb_loopi2_io_Out_2_ready = br_4_io_enable_ready; // @[bbgemm.scala 529:18]
  assign bb_loopi2_io_predicateIn_0_valid = Loop_3_io_activate_loop_start_valid; // @[bbgemm.scala 307:31]
  assign bb_loopi2_io_predicateIn_0_bits_taskID = Loop_3_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 307:31]
  assign bb_loopi2_io_predicateIn_0_bits_control = Loop_3_io_activate_loop_start_bits_control; // @[bbgemm.scala 307:31]
  assign bb_loopi2_io_predicateIn_1_valid = Loop_3_io_activate_loop_back_valid; // @[bbgemm.scala 309:31]
  assign bb_loopi2_io_predicateIn_1_bits_taskID = Loop_3_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 309:31]
  assign bb_loopi2_io_predicateIn_1_bits_control = Loop_3_io_activate_loop_back_bits_control; // @[bbgemm.scala 309:31]
  assign bb_loopk3_clock = clock;
  assign bb_loopk3_reset = reset;
  assign bb_loopk3_io_MaskBB_0_ready = phiindvars_iv785_io_Mask_ready; // @[bbgemm.scala 689:28]
  assign bb_loopk3_io_Out_0_ready = const2_io_enable_ready; // @[bbgemm.scala 532:20]
  assign bb_loopk3_io_Out_1_ready = const3_io_enable_ready; // @[bbgemm.scala 534:20]
  assign bb_loopk3_io_Out_2_ready = phiindvars_iv785_io_enable_ready; // @[bbgemm.scala 536:30]
  assign bb_loopk3_io_Out_3_ready = binaryOp_6_io_enable_ready; // @[bbgemm.scala 539:24]
  assign bb_loopk3_io_Out_4_ready = br_7_io_enable_ready; // @[bbgemm.scala 542:18]
  assign bb_loopk3_io_predicateIn_0_valid = Loop_2_io_activate_loop_back_valid; // @[bbgemm.scala 313:31]
  assign bb_loopk3_io_predicateIn_0_bits_taskID = Loop_2_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 313:31]
  assign bb_loopk3_io_predicateIn_0_bits_control = Loop_2_io_activate_loop_back_bits_control; // @[bbgemm.scala 313:31]
  assign bb_loopk3_io_predicateIn_1_valid = Loop_2_io_activate_loop_start_valid; // @[bbgemm.scala 311:31]
  assign bb_loopk3_io_predicateIn_1_bits_taskID = Loop_2_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 311:31]
  assign bb_loopk3_io_predicateIn_1_bits_control = Loop_2_io_activate_loop_start_bits_control; // @[bbgemm.scala 311:31]
  assign bb_for_body94_clock = clock;
  assign bb_for_body94_reset = reset;
  assign bb_for_body94_io_MaskBB_0_ready = phiindvars_iv718_io_Mask_ready; // @[bbgemm.scala 691:28]
  assign bb_for_body94_io_Out_0_ready = const4_io_enable_ready; // @[bbgemm.scala 545:20]
  assign bb_for_body94_io_Out_1_ready = const5_io_enable_ready; // @[bbgemm.scala 547:20]
  assign bb_for_body94_io_Out_2_ready = phiindvars_iv718_io_enable_ready; // @[bbgemm.scala 549:30]
  assign bb_for_body94_io_Out_3_ready = binaryOp_9_io_enable_ready; // @[bbgemm.scala 552:24]
  assign bb_for_body94_io_Out_4_ready = binaryOp_10_io_enable_ready; // @[bbgemm.scala 555:25]
  assign bb_for_body94_io_Out_5_ready = binaryOp_11_io_enable_ready; // @[bbgemm.scala 558:25]
  assign bb_for_body94_io_Out_6_ready = binaryOp_12_io_enable_ready; // @[bbgemm.scala 561:25]
  assign bb_for_body94_io_Out_7_ready = Gep_arrayidx13_io_enable_ready; // @[bbgemm.scala 564:28]
  assign bb_for_body94_io_Out_8_ready = ld_14_io_enable_ready; // @[bbgemm.scala 567:19]
  assign bb_for_body94_io_Out_9_ready = br_15_io_enable_ready; // @[bbgemm.scala 570:19]
  assign bb_for_body94_io_predicateIn_0_valid = Loop_1_io_activate_loop_back_valid; // @[bbgemm.scala 317:35]
  assign bb_for_body94_io_predicateIn_0_bits_taskID = Loop_1_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 317:35]
  assign bb_for_body94_io_predicateIn_0_bits_control = Loop_1_io_activate_loop_back_bits_control; // @[bbgemm.scala 317:35]
  assign bb_for_body94_io_predicateIn_1_valid = Loop_1_io_activate_loop_start_valid; // @[bbgemm.scala 315:35]
  assign bb_for_body94_io_predicateIn_1_bits_taskID = Loop_1_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 315:35]
  assign bb_for_body94_io_predicateIn_1_bits_control = Loop_1_io_activate_loop_start_bits_control; // @[bbgemm.scala 315:35]
  assign bb_for_body165_clock = clock;
  assign bb_for_body165_reset = reset;
  assign bb_for_body165_io_MaskBB_0_ready = phiindvars_iv16_io_Mask_ready; // @[bbgemm.scala 693:27]
  assign bb_for_body165_io_Out_0_ready = const6_io_enable_ready; // @[bbgemm.scala 573:20]
  assign bb_for_body165_io_Out_1_ready = const7_io_enable_ready; // @[bbgemm.scala 575:20]
  assign bb_for_body165_io_Out_2_ready = const8_io_enable_ready; // @[bbgemm.scala 577:20]
  assign bb_for_body165_io_Out_3_ready = phiindvars_iv16_io_enable_ready; // @[bbgemm.scala 579:29]
  assign bb_for_body165_io_Out_4_ready = binaryOp_17_io_enable_ready; // @[bbgemm.scala 582:25]
  assign bb_for_body165_io_Out_5_ready = binaryOp_18_io_enable_ready; // @[bbgemm.scala 585:25]
  assign bb_for_body165_io_Out_6_ready = Gep_arrayidx2019_io_enable_ready; // @[bbgemm.scala 588:30]
  assign bb_for_body165_io_Out_7_ready = ld_20_io_enable_ready; // @[bbgemm.scala 591:19]
  assign bb_for_body165_io_Out_8_ready = FP_mul2121_io_enable_ready; // @[bbgemm.scala 594:24]
  assign bb_for_body165_io_Out_9_ready = binaryOp_22_io_enable_ready; // @[bbgemm.scala 597:25]
  assign bb_for_body165_io_Out_10_ready = binaryOp_23_io_enable_ready; // @[bbgemm.scala 600:25]
  assign bb_for_body165_io_Out_11_ready = Gep_arrayidx2524_io_enable_ready; // @[bbgemm.scala 603:30]
  assign bb_for_body165_io_Out_12_ready = ld_25_io_enable_ready; // @[bbgemm.scala 606:19]
  assign bb_for_body165_io_Out_13_ready = FP_add2626_io_enable_ready; // @[bbgemm.scala 609:24]
  assign bb_for_body165_io_Out_14_ready = st_27_io_enable_ready; // @[bbgemm.scala 612:19]
  assign bb_for_body165_io_Out_15_ready = binaryOp_indvars_iv_next28_io_enable_ready; // @[bbgemm.scala 615:40]
  assign bb_for_body165_io_Out_16_ready = icmp_exitcond29_io_enable_ready; // @[bbgemm.scala 618:29]
  assign bb_for_body165_io_Out_17_ready = br_30_io_enable_ready; // @[bbgemm.scala 621:19]
  assign bb_for_body165_io_predicateIn_0_valid = Loop_0_io_activate_loop_back_valid; // @[bbgemm.scala 321:36]
  assign bb_for_body165_io_predicateIn_0_bits_taskID = Loop_0_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 321:36]
  assign bb_for_body165_io_predicateIn_0_bits_control = Loop_0_io_activate_loop_back_bits_control; // @[bbgemm.scala 321:36]
  assign bb_for_body165_io_predicateIn_1_valid = Loop_0_io_activate_loop_start_valid; // @[bbgemm.scala 319:36]
  assign bb_for_body165_io_predicateIn_1_bits_taskID = Loop_0_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 319:36]
  assign bb_for_body165_io_predicateIn_1_bits_control = Loop_0_io_activate_loop_start_bits_control; // @[bbgemm.scala 319:36]
  assign bb_for_inc276_clock = clock;
  assign bb_for_inc276_reset = reset;
  assign bb_for_inc276_io_predicateIn_0_valid = Loop_0_io_loopExit_0_valid; // @[bbgemm.scala 323:35]
  assign bb_for_inc276_io_predicateIn_0_bits_taskID = Loop_0_io_loopExit_0_bits_taskID; // @[bbgemm.scala 323:35]
  assign bb_for_inc276_io_predicateIn_0_bits_control = Loop_0_io_loopExit_0_bits_control; // @[bbgemm.scala 323:35]
  assign bb_for_inc276_io_Out_0_ready = const9_io_enable_ready; // @[bbgemm.scala 624:20]
  assign bb_for_inc276_io_Out_1_ready = const10_io_enable_ready; // @[bbgemm.scala 626:21]
  assign bb_for_inc276_io_Out_2_ready = binaryOp_indvars_iv_next7231_io_enable_ready; // @[bbgemm.scala 628:42]
  assign bb_for_inc276_io_Out_3_ready = icmp_exitcond7732_io_enable_ready; // @[bbgemm.scala 631:31]
  assign bb_for_inc276_io_Out_4_ready = br_33_io_enable_ready; // @[bbgemm.scala 634:19]
  assign bb_for_inc307_clock = clock;
  assign bb_for_inc307_reset = reset;
  assign bb_for_inc307_io_predicateIn_0_valid = Loop_1_io_loopExit_0_valid; // @[bbgemm.scala 325:35]
  assign bb_for_inc307_io_predicateIn_0_bits_taskID = Loop_1_io_loopExit_0_bits_taskID; // @[bbgemm.scala 325:35]
  assign bb_for_inc307_io_predicateIn_0_bits_control = Loop_1_io_loopExit_0_bits_control; // @[bbgemm.scala 325:35]
  assign bb_for_inc307_io_Out_0_ready = const11_io_enable_ready; // @[bbgemm.scala 637:21]
  assign bb_for_inc307_io_Out_1_ready = const12_io_enable_ready; // @[bbgemm.scala 639:21]
  assign bb_for_inc307_io_Out_2_ready = binaryOp_indvars_iv_next7934_io_enable_ready; // @[bbgemm.scala 641:42]
  assign bb_for_inc307_io_Out_3_ready = icmp_exitcond8135_io_enable_ready; // @[bbgemm.scala 644:31]
  assign bb_for_inc307_io_Out_4_ready = br_36_io_enable_ready; // @[bbgemm.scala 647:19]
  assign bb_for_inc338_clock = clock;
  assign bb_for_inc338_reset = reset;
  assign bb_for_inc338_io_predicateIn_0_valid = Loop_2_io_loopExit_0_valid; // @[bbgemm.scala 327:35]
  assign bb_for_inc338_io_predicateIn_0_bits_taskID = Loop_2_io_loopExit_0_bits_taskID; // @[bbgemm.scala 327:35]
  assign bb_for_inc338_io_predicateIn_0_bits_control = Loop_2_io_loopExit_0_bits_control; // @[bbgemm.scala 327:35]
  assign bb_for_inc338_io_Out_0_ready = const13_io_enable_ready; // @[bbgemm.scala 650:21]
  assign bb_for_inc338_io_Out_1_ready = const14_io_enable_ready; // @[bbgemm.scala 652:21]
  assign bb_for_inc338_io_Out_2_ready = binaryOp_indvars_iv_next8337_io_enable_ready; // @[bbgemm.scala 654:42]
  assign bb_for_inc338_io_Out_3_ready = icmp_cmp238_io_enable_ready; // @[bbgemm.scala 657:25]
  assign bb_for_inc338_io_Out_4_ready = br_39_io_enable_ready; // @[bbgemm.scala 660:19]
  assign bb_for_inc369_clock = clock;
  assign bb_for_inc369_reset = reset;
  assign bb_for_inc369_io_predicateIn_0_valid = Loop_3_io_loopExit_0_valid; // @[bbgemm.scala 329:35]
  assign bb_for_inc369_io_predicateIn_0_bits_taskID = Loop_3_io_loopExit_0_bits_taskID; // @[bbgemm.scala 329:35]
  assign bb_for_inc369_io_predicateIn_0_bits_control = Loop_3_io_loopExit_0_bits_control; // @[bbgemm.scala 329:35]
  assign bb_for_inc369_io_Out_0_ready = const15_io_enable_ready; // @[bbgemm.scala 663:21]
  assign bb_for_inc369_io_Out_1_ready = const16_io_enable_ready; // @[bbgemm.scala 665:21]
  assign bb_for_inc369_io_Out_2_ready = binaryOp_indvars_iv_next8540_io_enable_ready; // @[bbgemm.scala 667:42]
  assign bb_for_inc369_io_Out_3_ready = icmp_cmp41_io_enable_ready; // @[bbgemm.scala 670:24]
  assign bb_for_inc369_io_Out_4_ready = br_42_io_enable_ready; // @[bbgemm.scala 673:19]
  assign bb_for_end3810_clock = clock;
  assign bb_for_end3810_reset = reset;
  assign bb_for_end3810_io_predicateIn_0_valid = Loop_4_io_loopExit_0_valid; // @[bbgemm.scala 331:36]
  assign bb_for_end3810_io_predicateIn_0_bits_taskID = Loop_4_io_loopExit_0_bits_taskID; // @[bbgemm.scala 331:36]
  assign bb_for_end3810_io_predicateIn_0_bits_control = Loop_4_io_loopExit_0_bits_control; // @[bbgemm.scala 331:36]
  assign bb_for_end3810_io_Out_0_ready = ret_43_io_In_enable_ready; // @[bbgemm.scala 676:23]
  assign br_0_clock = clock;
  assign br_0_reset = reset;
  assign br_0_io_enable_valid = bb_entry0_io_Out_0_valid; // @[bbgemm.scala 513:18]
  assign br_0_io_enable_bits_control = bb_entry0_io_Out_0_bits_control; // @[bbgemm.scala 513:18]
  assign br_0_io_Out_0_ready = Loop_4_io_enable_ready; // @[bbgemm.scala 369:20]
  assign phiindvars_iv841_clock = clock;
  assign phiindvars_iv841_reset = reset;
  assign phiindvars_iv841_io_enable_valid = bb_loopkk1_io_Out_1_valid; // @[bbgemm.scala 518:30]
  assign phiindvars_iv841_io_enable_bits_control = bb_loopkk1_io_Out_1_bits_control; // @[bbgemm.scala 518:30]
  assign phiindvars_iv841_io_InData_0_valid = const0_io_Out_valid; // @[bbgemm.scala 734:33]
  assign phiindvars_iv841_io_InData_0_bits_taskID = const0_io_Out_bits_taskID; // @[bbgemm.scala 734:33]
  assign phiindvars_iv841_io_InData_1_valid = Loop_4_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 505:33]
  assign phiindvars_iv841_io_InData_1_bits_taskID = Loop_4_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 505:33]
  assign phiindvars_iv841_io_InData_1_bits_data = Loop_4_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 505:33]
  assign phiindvars_iv841_io_Mask_valid = bb_loopkk1_io_MaskBB_0_valid; // @[bbgemm.scala 685:28]
  assign phiindvars_iv841_io_Mask_bits = bb_loopkk1_io_MaskBB_0_bits; // @[bbgemm.scala 685:28]
  assign phiindvars_iv841_io_Out_0_ready = Loop_3_io_InLiveIn_0_ready; // @[bbgemm.scala 421:25]
  assign phiindvars_iv841_io_Out_1_ready = binaryOp_indvars_iv_next8540_io_LeftIO_ready; // @[bbgemm.scala 768:42]
  assign br_2_clock = clock;
  assign br_2_reset = reset;
  assign br_2_io_enable_valid = bb_loopkk1_io_Out_2_valid; // @[bbgemm.scala 521:18]
  assign br_2_io_enable_bits_taskID = bb_loopkk1_io_Out_2_bits_taskID; // @[bbgemm.scala 521:18]
  assign br_2_io_enable_bits_control = bb_loopkk1_io_Out_2_bits_control; // @[bbgemm.scala 521:18]
  assign br_2_io_Out_0_ready = Loop_3_io_enable_ready; // @[bbgemm.scala 363:20]
  assign phiindvars_iv823_clock = clock;
  assign phiindvars_iv823_reset = reset;
  assign phiindvars_iv823_io_enable_valid = bb_loopi2_io_Out_1_valid; // @[bbgemm.scala 526:30]
  assign phiindvars_iv823_io_enable_bits_control = bb_loopi2_io_Out_1_bits_control; // @[bbgemm.scala 526:30]
  assign phiindvars_iv823_io_InData_0_valid = const1_io_Out_valid; // @[bbgemm.scala 736:33]
  assign phiindvars_iv823_io_InData_0_bits_taskID = const1_io_Out_bits_taskID; // @[bbgemm.scala 736:33]
  assign phiindvars_iv823_io_InData_1_valid = Loop_3_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 503:33]
  assign phiindvars_iv823_io_InData_1_bits_taskID = Loop_3_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 503:33]
  assign phiindvars_iv823_io_InData_1_bits_data = Loop_3_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 503:33]
  assign phiindvars_iv823_io_Mask_valid = bb_loopi2_io_MaskBB_0_valid; // @[bbgemm.scala 687:28]
  assign phiindvars_iv823_io_Mask_bits = bb_loopi2_io_MaskBB_0_bits; // @[bbgemm.scala 687:28]
  assign phiindvars_iv823_io_Out_0_ready = Loop_2_io_InLiveIn_0_ready; // @[bbgemm.scala 411:25]
  assign phiindvars_iv823_io_Out_1_ready = binaryOp_indvars_iv_next8337_io_LeftIO_ready; // @[bbgemm.scala 770:42]
  assign br_4_clock = clock;
  assign br_4_reset = reset;
  assign br_4_io_enable_valid = bb_loopi2_io_Out_2_valid; // @[bbgemm.scala 529:18]
  assign br_4_io_enable_bits_taskID = bb_loopi2_io_Out_2_bits_taskID; // @[bbgemm.scala 529:18]
  assign br_4_io_enable_bits_control = bb_loopi2_io_Out_2_bits_control; // @[bbgemm.scala 529:18]
  assign br_4_io_Out_0_ready = Loop_2_io_enable_ready; // @[bbgemm.scala 357:20]
  assign phiindvars_iv785_clock = clock;
  assign phiindvars_iv785_reset = reset;
  assign phiindvars_iv785_io_enable_valid = bb_loopk3_io_Out_2_valid; // @[bbgemm.scala 536:30]
  assign phiindvars_iv785_io_enable_bits_control = bb_loopk3_io_Out_2_bits_control; // @[bbgemm.scala 536:30]
  assign phiindvars_iv785_io_InData_0_valid = const2_io_Out_valid; // @[bbgemm.scala 738:33]
  assign phiindvars_iv785_io_InData_0_bits_taskID = const2_io_Out_bits_taskID; // @[bbgemm.scala 738:33]
  assign phiindvars_iv785_io_InData_1_valid = Loop_2_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 501:33]
  assign phiindvars_iv785_io_InData_1_bits_taskID = Loop_2_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 501:33]
  assign phiindvars_iv785_io_InData_1_bits_data = Loop_2_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 501:33]
  assign phiindvars_iv785_io_Mask_valid = bb_loopk3_io_MaskBB_0_valid; // @[bbgemm.scala 689:28]
  assign phiindvars_iv785_io_Mask_bits = bb_loopk3_io_MaskBB_0_bits; // @[bbgemm.scala 689:28]
  assign phiindvars_iv785_io_Out_0_ready = binaryOp_6_io_LeftIO_ready; // @[bbgemm.scala 772:24]
  assign phiindvars_iv785_io_Out_1_ready = binaryOp_indvars_iv_next7934_io_LeftIO_ready; // @[bbgemm.scala 774:42]
  assign binaryOp_6_clock = clock;
  assign binaryOp_6_reset = reset;
  assign binaryOp_6_io_enable_valid = bb_loopk3_io_Out_3_valid; // @[bbgemm.scala 539:24]
  assign binaryOp_6_io_enable_bits_taskID = bb_loopk3_io_Out_3_bits_taskID; // @[bbgemm.scala 539:24]
  assign binaryOp_6_io_enable_bits_control = bb_loopk3_io_Out_3_bits_control; // @[bbgemm.scala 539:24]
  assign binaryOp_6_io_Out_0_ready = Loop_1_io_InLiveIn_0_ready; // @[bbgemm.scala 399:25]
  assign binaryOp_6_io_LeftIO_valid = phiindvars_iv785_io_Out_0_valid; // @[bbgemm.scala 772:24]
  assign binaryOp_6_io_LeftIO_bits_data = phiindvars_iv785_io_Out_0_bits_data; // @[bbgemm.scala 772:24]
  assign binaryOp_6_io_RightIO_valid = const3_io_Out_valid; // @[bbgemm.scala 740:25]
  assign br_7_clock = clock;
  assign br_7_reset = reset;
  assign br_7_io_enable_valid = bb_loopk3_io_Out_4_valid; // @[bbgemm.scala 542:18]
  assign br_7_io_enable_bits_taskID = bb_loopk3_io_Out_4_bits_taskID; // @[bbgemm.scala 542:18]
  assign br_7_io_enable_bits_control = bb_loopk3_io_Out_4_bits_control; // @[bbgemm.scala 542:18]
  assign br_7_io_Out_0_ready = Loop_1_io_enable_ready; // @[bbgemm.scala 351:20]
  assign phiindvars_iv718_clock = clock;
  assign phiindvars_iv718_reset = reset;
  assign phiindvars_iv718_io_enable_valid = bb_for_body94_io_Out_2_valid; // @[bbgemm.scala 549:30]
  assign phiindvars_iv718_io_enable_bits_control = bb_for_body94_io_Out_2_bits_control; // @[bbgemm.scala 549:30]
  assign phiindvars_iv718_io_InData_0_valid = const4_io_Out_valid; // @[bbgemm.scala 742:33]
  assign phiindvars_iv718_io_InData_0_bits_taskID = const4_io_Out_bits_taskID; // @[bbgemm.scala 742:33]
  assign phiindvars_iv718_io_InData_1_valid = Loop_1_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 499:33]
  assign phiindvars_iv718_io_InData_1_bits_taskID = Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 499:33]
  assign phiindvars_iv718_io_InData_1_bits_data = Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 499:33]
  assign phiindvars_iv718_io_Mask_valid = bb_for_body94_io_MaskBB_0_valid; // @[bbgemm.scala 691:28]
  assign phiindvars_iv718_io_Mask_bits = bb_for_body94_io_MaskBB_0_bits; // @[bbgemm.scala 691:28]
  assign phiindvars_iv718_io_Out_0_ready = binaryOp_9_io_LeftIO_ready; // @[bbgemm.scala 776:24]
  assign phiindvars_iv718_io_Out_1_ready = binaryOp_11_io_LeftIO_ready; // @[bbgemm.scala 778:25]
  assign phiindvars_iv718_io_Out_2_ready = binaryOp_indvars_iv_next7231_io_LeftIO_ready; // @[bbgemm.scala 780:42]
  assign binaryOp_9_clock = clock;
  assign binaryOp_9_reset = reset;
  assign binaryOp_9_io_enable_valid = bb_for_body94_io_Out_3_valid; // @[bbgemm.scala 552:24]
  assign binaryOp_9_io_enable_bits_taskID = bb_for_body94_io_Out_3_bits_taskID; // @[bbgemm.scala 552:24]
  assign binaryOp_9_io_enable_bits_control = bb_for_body94_io_Out_3_bits_control; // @[bbgemm.scala 552:24]
  assign binaryOp_9_io_Out_0_ready = binaryOp_10_io_LeftIO_ready; // @[bbgemm.scala 782:25]
  assign binaryOp_9_io_LeftIO_valid = phiindvars_iv718_io_Out_0_valid; // @[bbgemm.scala 776:24]
  assign binaryOp_9_io_LeftIO_bits_data = phiindvars_iv718_io_Out_0_bits_data; // @[bbgemm.scala 776:24]
  assign binaryOp_9_io_RightIO_valid = Loop_1_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 457:25]
  assign binaryOp_9_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 457:25]
  assign binaryOp_10_clock = clock;
  assign binaryOp_10_reset = reset;
  assign binaryOp_10_io_enable_valid = bb_for_body94_io_Out_4_valid; // @[bbgemm.scala 555:25]
  assign binaryOp_10_io_enable_bits_taskID = bb_for_body94_io_Out_4_bits_taskID; // @[bbgemm.scala 555:25]
  assign binaryOp_10_io_enable_bits_control = bb_for_body94_io_Out_4_bits_control; // @[bbgemm.scala 555:25]
  assign binaryOp_10_io_Out_0_ready = Loop_0_io_InLiveIn_0_ready; // @[bbgemm.scala 387:25]
  assign binaryOp_10_io_LeftIO_valid = binaryOp_9_io_Out_0_valid; // @[bbgemm.scala 782:25]
  assign binaryOp_10_io_LeftIO_bits_data = binaryOp_9_io_Out_0_bits_data; // @[bbgemm.scala 782:25]
  assign binaryOp_10_io_RightIO_valid = const5_io_Out_valid; // @[bbgemm.scala 744:26]
  assign binaryOp_11_clock = clock;
  assign binaryOp_11_reset = reset;
  assign binaryOp_11_io_enable_valid = bb_for_body94_io_Out_5_valid; // @[bbgemm.scala 558:25]
  assign binaryOp_11_io_enable_bits_taskID = bb_for_body94_io_Out_5_bits_taskID; // @[bbgemm.scala 558:25]
  assign binaryOp_11_io_enable_bits_control = bb_for_body94_io_Out_5_bits_control; // @[bbgemm.scala 558:25]
  assign binaryOp_11_io_Out_0_ready = binaryOp_12_io_LeftIO_ready; // @[bbgemm.scala 784:25]
  assign binaryOp_11_io_LeftIO_valid = phiindvars_iv718_io_Out_1_valid; // @[bbgemm.scala 778:25]
  assign binaryOp_11_io_LeftIO_bits_data = phiindvars_iv718_io_Out_1_bits_data; // @[bbgemm.scala 778:25]
  assign binaryOp_11_io_RightIO_valid = Loop_1_io_OutLiveIn_field4_1_valid; // @[bbgemm.scala 459:26]
  assign binaryOp_11_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field4_1_bits_data; // @[bbgemm.scala 459:26]
  assign binaryOp_12_clock = clock;
  assign binaryOp_12_reset = reset;
  assign binaryOp_12_io_enable_valid = bb_for_body94_io_Out_6_valid; // @[bbgemm.scala 561:25]
  assign binaryOp_12_io_enable_bits_taskID = bb_for_body94_io_Out_6_bits_taskID; // @[bbgemm.scala 561:25]
  assign binaryOp_12_io_enable_bits_control = bb_for_body94_io_Out_6_bits_control; // @[bbgemm.scala 561:25]
  assign binaryOp_12_io_Out_0_ready = Gep_arrayidx13_io_idx_0_ready; // @[bbgemm.scala 786:28]
  assign binaryOp_12_io_LeftIO_valid = binaryOp_11_io_Out_0_valid; // @[bbgemm.scala 784:25]
  assign binaryOp_12_io_LeftIO_bits_data = binaryOp_11_io_Out_0_bits_data; // @[bbgemm.scala 784:25]
  assign binaryOp_12_io_RightIO_valid = Loop_1_io_OutLiveIn_field0_1_valid; // @[bbgemm.scala 455:26]
  assign binaryOp_12_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field0_1_bits_data; // @[bbgemm.scala 455:26]
  assign Gep_arrayidx13_clock = clock;
  assign Gep_arrayidx13_reset = reset;
  assign Gep_arrayidx13_io_enable_valid = bb_for_body94_io_Out_7_valid; // @[bbgemm.scala 564:28]
  assign Gep_arrayidx13_io_enable_bits_taskID = bb_for_body94_io_Out_7_bits_taskID; // @[bbgemm.scala 564:28]
  assign Gep_arrayidx13_io_enable_bits_control = bb_for_body94_io_Out_7_bits_control; // @[bbgemm.scala 564:28]
  assign Gep_arrayidx13_io_Out_0_ready = ld_14_io_GepAddr_ready; // @[bbgemm.scala 788:20]
  assign Gep_arrayidx13_io_baseAddress_valid = Loop_1_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 461:33]
  assign Gep_arrayidx13_io_baseAddress_bits_data = Loop_1_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 461:33]
  assign Gep_arrayidx13_io_idx_0_valid = binaryOp_12_io_Out_0_valid; // @[bbgemm.scala 786:28]
  assign Gep_arrayidx13_io_idx_0_bits_data = binaryOp_12_io_Out_0_bits_data; // @[bbgemm.scala 786:28]
  assign ld_14_clock = clock;
  assign ld_14_reset = reset;
  assign ld_14_io_enable_valid = bb_for_body94_io_Out_8_valid; // @[bbgemm.scala 567:19]
  assign ld_14_io_enable_bits_taskID = bb_for_body94_io_Out_8_bits_taskID; // @[bbgemm.scala 567:19]
  assign ld_14_io_enable_bits_control = bb_for_body94_io_Out_8_bits_control; // @[bbgemm.scala 567:19]
  assign ld_14_io_Out_0_ready = Loop_0_io_InLiveIn_1_ready; // @[bbgemm.scala 389:25]
  assign ld_14_io_GepAddr_valid = Gep_arrayidx13_io_Out_0_valid; // @[bbgemm.scala 788:20]
  assign ld_14_io_GepAddr_bits_data = Gep_arrayidx13_io_Out_0_bits_data; // @[bbgemm.scala 788:20]
  assign ld_14_io_MemReq_ready = MemCtrl_io_rd_mem_0_MemReq_ready; // @[bbgemm.scala 707:31]
  assign ld_14_io_MemResp_valid = MemCtrl_io_rd_mem_0_MemResp_valid; // @[bbgemm.scala 709:20]
  assign ld_14_io_MemResp_bits_data = MemCtrl_io_rd_mem_0_MemResp_bits_data; // @[bbgemm.scala 709:20]
  assign br_15_clock = clock;
  assign br_15_reset = reset;
  assign br_15_io_enable_valid = bb_for_body94_io_Out_9_valid; // @[bbgemm.scala 570:19]
  assign br_15_io_enable_bits_taskID = bb_for_body94_io_Out_9_bits_taskID; // @[bbgemm.scala 570:19]
  assign br_15_io_enable_bits_control = bb_for_body94_io_Out_9_bits_control; // @[bbgemm.scala 570:19]
  assign br_15_io_Out_0_ready = Loop_0_io_enable_ready; // @[bbgemm.scala 345:20]
  assign phiindvars_iv16_clock = clock;
  assign phiindvars_iv16_reset = reset;
  assign phiindvars_iv16_io_enable_valid = bb_for_body165_io_Out_3_valid; // @[bbgemm.scala 579:29]
  assign phiindvars_iv16_io_enable_bits_control = bb_for_body165_io_Out_3_bits_control; // @[bbgemm.scala 579:29]
  assign phiindvars_iv16_io_InData_0_valid = const6_io_Out_valid; // @[bbgemm.scala 746:32]
  assign phiindvars_iv16_io_InData_0_bits_taskID = const6_io_Out_bits_taskID; // @[bbgemm.scala 746:32]
  assign phiindvars_iv16_io_InData_1_valid = Loop_0_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 497:32]
  assign phiindvars_iv16_io_InData_1_bits_taskID = Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 497:32]
  assign phiindvars_iv16_io_InData_1_bits_data = Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 497:32]
  assign phiindvars_iv16_io_Mask_valid = bb_for_body165_io_MaskBB_0_valid; // @[bbgemm.scala 693:27]
  assign phiindvars_iv16_io_Mask_bits = bb_for_body165_io_MaskBB_0_bits; // @[bbgemm.scala 693:27]
  assign phiindvars_iv16_io_Out_0_ready = binaryOp_17_io_LeftIO_ready; // @[bbgemm.scala 790:25]
  assign phiindvars_iv16_io_Out_1_ready = binaryOp_22_io_LeftIO_ready; // @[bbgemm.scala 792:25]
  assign phiindvars_iv16_io_Out_2_ready = binaryOp_indvars_iv_next28_io_LeftIO_ready; // @[bbgemm.scala 794:40]
  assign binaryOp_17_clock = clock;
  assign binaryOp_17_reset = reset;
  assign binaryOp_17_io_enable_valid = bb_for_body165_io_Out_4_valid; // @[bbgemm.scala 582:25]
  assign binaryOp_17_io_enable_bits_taskID = bb_for_body165_io_Out_4_bits_taskID; // @[bbgemm.scala 582:25]
  assign binaryOp_17_io_enable_bits_control = bb_for_body165_io_Out_4_bits_control; // @[bbgemm.scala 582:25]
  assign binaryOp_17_io_Out_0_ready = binaryOp_18_io_LeftIO_ready; // @[bbgemm.scala 796:25]
  assign binaryOp_17_io_LeftIO_valid = phiindvars_iv16_io_Out_0_valid; // @[bbgemm.scala 790:25]
  assign binaryOp_17_io_LeftIO_bits_data = phiindvars_iv16_io_Out_0_bits_data; // @[bbgemm.scala 790:25]
  assign binaryOp_17_io_RightIO_valid = Loop_0_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 451:26]
  assign binaryOp_17_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 451:26]
  assign binaryOp_18_clock = clock;
  assign binaryOp_18_reset = reset;
  assign binaryOp_18_io_enable_valid = bb_for_body165_io_Out_5_valid; // @[bbgemm.scala 585:25]
  assign binaryOp_18_io_enable_bits_taskID = bb_for_body165_io_Out_5_bits_taskID; // @[bbgemm.scala 585:25]
  assign binaryOp_18_io_enable_bits_control = bb_for_body165_io_Out_5_bits_control; // @[bbgemm.scala 585:25]
  assign binaryOp_18_io_Out_0_ready = Gep_arrayidx2019_io_idx_0_ready; // @[bbgemm.scala 798:30]
  assign binaryOp_18_io_LeftIO_valid = binaryOp_17_io_Out_0_valid; // @[bbgemm.scala 796:25]
  assign binaryOp_18_io_LeftIO_bits_data = binaryOp_17_io_Out_0_bits_data; // @[bbgemm.scala 796:25]
  assign binaryOp_18_io_RightIO_valid = Loop_0_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 441:26]
  assign binaryOp_18_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 441:26]
  assign Gep_arrayidx2019_clock = clock;
  assign Gep_arrayidx2019_reset = reset;
  assign Gep_arrayidx2019_io_enable_valid = bb_for_body165_io_Out_6_valid; // @[bbgemm.scala 588:30]
  assign Gep_arrayidx2019_io_enable_bits_taskID = bb_for_body165_io_Out_6_bits_taskID; // @[bbgemm.scala 588:30]
  assign Gep_arrayidx2019_io_enable_bits_control = bb_for_body165_io_Out_6_bits_control; // @[bbgemm.scala 588:30]
  assign Gep_arrayidx2019_io_Out_0_ready = ld_20_io_GepAddr_ready; // @[bbgemm.scala 800:20]
  assign Gep_arrayidx2019_io_baseAddress_valid = Loop_0_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 445:35]
  assign Gep_arrayidx2019_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 445:35]
  assign Gep_arrayidx2019_io_idx_0_valid = binaryOp_18_io_Out_0_valid; // @[bbgemm.scala 798:30]
  assign Gep_arrayidx2019_io_idx_0_bits_data = binaryOp_18_io_Out_0_bits_data; // @[bbgemm.scala 798:30]
  assign ld_20_clock = clock;
  assign ld_20_reset = reset;
  assign ld_20_io_enable_valid = bb_for_body165_io_Out_7_valid; // @[bbgemm.scala 591:19]
  assign ld_20_io_enable_bits_taskID = bb_for_body165_io_Out_7_bits_taskID; // @[bbgemm.scala 591:19]
  assign ld_20_io_enable_bits_control = bb_for_body165_io_Out_7_bits_control; // @[bbgemm.scala 591:19]
  assign ld_20_io_Out_0_ready = FP_mul2121_io_RightIO_ready; // @[bbgemm.scala 802:25]
  assign ld_20_io_GepAddr_valid = Gep_arrayidx2019_io_Out_0_valid; // @[bbgemm.scala 800:20]
  assign ld_20_io_GepAddr_bits_data = Gep_arrayidx2019_io_Out_0_bits_data; // @[bbgemm.scala 800:20]
  assign ld_20_io_MemReq_ready = MemCtrl_io_rd_mem_1_MemReq_ready; // @[bbgemm.scala 711:31]
  assign ld_20_io_MemResp_valid = MemCtrl_io_rd_mem_1_MemResp_valid; // @[bbgemm.scala 713:20]
  assign ld_20_io_MemResp_bits_data = MemCtrl_io_rd_mem_1_MemResp_bits_data; // @[bbgemm.scala 713:20]
  assign FP_mul2121_clock = clock;
  assign FP_mul2121_reset = reset;
  assign FP_mul2121_io_enable_valid = bb_for_body165_io_Out_8_valid; // @[bbgemm.scala 594:24]
  assign FP_mul2121_io_enable_bits_taskID = bb_for_body165_io_Out_8_bits_taskID; // @[bbgemm.scala 594:24]
  assign FP_mul2121_io_enable_bits_control = bb_for_body165_io_Out_8_bits_control; // @[bbgemm.scala 594:24]
  assign FP_mul2121_io_Out_0_ready = FP_add2626_io_RightIO_ready; // @[bbgemm.scala 804:25]
  assign FP_mul2121_io_LeftIO_valid = Loop_0_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 443:24]
  assign FP_mul2121_io_LeftIO_bits_data = Loop_0_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 443:24]
  assign FP_mul2121_io_RightIO_valid = ld_20_io_Out_0_valid; // @[bbgemm.scala 802:25]
  assign FP_mul2121_io_RightIO_bits_data = ld_20_io_Out_0_bits_data; // @[bbgemm.scala 802:25]
  assign binaryOp_22_clock = clock;
  assign binaryOp_22_reset = reset;
  assign binaryOp_22_io_enable_valid = bb_for_body165_io_Out_9_valid; // @[bbgemm.scala 597:25]
  assign binaryOp_22_io_enable_bits_taskID = bb_for_body165_io_Out_9_bits_taskID; // @[bbgemm.scala 597:25]
  assign binaryOp_22_io_enable_bits_control = bb_for_body165_io_Out_9_bits_control; // @[bbgemm.scala 597:25]
  assign binaryOp_22_io_Out_0_ready = binaryOp_23_io_LeftIO_ready; // @[bbgemm.scala 806:25]
  assign binaryOp_22_io_LeftIO_valid = phiindvars_iv16_io_Out_1_valid; // @[bbgemm.scala 792:25]
  assign binaryOp_22_io_LeftIO_bits_data = phiindvars_iv16_io_Out_1_bits_data; // @[bbgemm.scala 792:25]
  assign binaryOp_22_io_RightIO_valid = Loop_0_io_OutLiveIn_field5_1_valid; // @[bbgemm.scala 453:26]
  assign binaryOp_22_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field5_1_bits_data; // @[bbgemm.scala 453:26]
  assign binaryOp_23_clock = clock;
  assign binaryOp_23_reset = reset;
  assign binaryOp_23_io_enable_valid = bb_for_body165_io_Out_10_valid; // @[bbgemm.scala 600:25]
  assign binaryOp_23_io_enable_bits_taskID = bb_for_body165_io_Out_10_bits_taskID; // @[bbgemm.scala 600:25]
  assign binaryOp_23_io_enable_bits_control = bb_for_body165_io_Out_10_bits_control; // @[bbgemm.scala 600:25]
  assign binaryOp_23_io_Out_0_ready = Gep_arrayidx2524_io_idx_0_ready; // @[bbgemm.scala 808:30]
  assign binaryOp_23_io_LeftIO_valid = binaryOp_22_io_Out_0_valid; // @[bbgemm.scala 806:25]
  assign binaryOp_23_io_LeftIO_bits_data = binaryOp_22_io_Out_0_bits_data; // @[bbgemm.scala 806:25]
  assign binaryOp_23_io_RightIO_valid = Loop_0_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 447:26]
  assign binaryOp_23_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 447:26]
  assign Gep_arrayidx2524_clock = clock;
  assign Gep_arrayidx2524_reset = reset;
  assign Gep_arrayidx2524_io_enable_valid = bb_for_body165_io_Out_11_valid; // @[bbgemm.scala 603:30]
  assign Gep_arrayidx2524_io_enable_bits_taskID = bb_for_body165_io_Out_11_bits_taskID; // @[bbgemm.scala 603:30]
  assign Gep_arrayidx2524_io_enable_bits_control = bb_for_body165_io_Out_11_bits_control; // @[bbgemm.scala 603:30]
  assign Gep_arrayidx2524_io_Out_0_ready = ld_25_io_GepAddr_ready; // @[bbgemm.scala 810:20]
  assign Gep_arrayidx2524_io_Out_1_ready = st_27_io_GepAddr_ready; // @[bbgemm.scala 812:20]
  assign Gep_arrayidx2524_io_baseAddress_valid = Loop_0_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 449:35]
  assign Gep_arrayidx2524_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 449:35]
  assign Gep_arrayidx2524_io_idx_0_valid = binaryOp_23_io_Out_0_valid; // @[bbgemm.scala 808:30]
  assign Gep_arrayidx2524_io_idx_0_bits_data = binaryOp_23_io_Out_0_bits_data; // @[bbgemm.scala 808:30]
  assign ld_25_clock = clock;
  assign ld_25_reset = reset;
  assign ld_25_io_enable_valid = bb_for_body165_io_Out_12_valid; // @[bbgemm.scala 606:19]
  assign ld_25_io_enable_bits_taskID = bb_for_body165_io_Out_12_bits_taskID; // @[bbgemm.scala 606:19]
  assign ld_25_io_enable_bits_control = bb_for_body165_io_Out_12_bits_control; // @[bbgemm.scala 606:19]
  assign ld_25_io_Out_0_ready = FP_add2626_io_LeftIO_ready; // @[bbgemm.scala 814:24]
  assign ld_25_io_GepAddr_valid = Gep_arrayidx2524_io_Out_0_valid; // @[bbgemm.scala 810:20]
  assign ld_25_io_GepAddr_bits_data = Gep_arrayidx2524_io_Out_0_bits_data; // @[bbgemm.scala 810:20]
  assign ld_25_io_MemReq_ready = MemCtrl_io_rd_mem_2_MemReq_ready; // @[bbgemm.scala 715:31]
  assign ld_25_io_MemResp_valid = MemCtrl_io_rd_mem_2_MemResp_valid; // @[bbgemm.scala 717:20]
  assign ld_25_io_MemResp_bits_data = MemCtrl_io_rd_mem_2_MemResp_bits_data; // @[bbgemm.scala 717:20]
  assign FP_add2626_clock = clock;
  assign FP_add2626_reset = reset;
  assign FP_add2626_io_enable_valid = bb_for_body165_io_Out_13_valid; // @[bbgemm.scala 609:24]
  assign FP_add2626_io_enable_bits_taskID = bb_for_body165_io_Out_13_bits_taskID; // @[bbgemm.scala 609:24]
  assign FP_add2626_io_enable_bits_control = bb_for_body165_io_Out_13_bits_control; // @[bbgemm.scala 609:24]
  assign FP_add2626_io_Out_0_ready = st_27_io_inData_ready; // @[bbgemm.scala 816:19]
  assign FP_add2626_io_LeftIO_valid = ld_25_io_Out_0_valid; // @[bbgemm.scala 814:24]
  assign FP_add2626_io_LeftIO_bits_data = ld_25_io_Out_0_bits_data; // @[bbgemm.scala 814:24]
  assign FP_add2626_io_RightIO_valid = FP_mul2121_io_Out_0_valid; // @[bbgemm.scala 804:25]
  assign FP_add2626_io_RightIO_bits_data = FP_mul2121_io_Out_0_bits_data; // @[bbgemm.scala 804:25]
  assign st_27_clock = clock;
  assign st_27_reset = reset;
  assign st_27_io_enable_valid = bb_for_body165_io_Out_14_valid; // @[bbgemm.scala 612:19]
  assign st_27_io_enable_bits_taskID = bb_for_body165_io_Out_14_bits_taskID; // @[bbgemm.scala 612:19]
  assign st_27_io_enable_bits_control = bb_for_body165_io_Out_14_bits_control; // @[bbgemm.scala 612:19]
  assign st_27_io_SuccOp_0_ready = br_30_io_PredOp_0_ready; // @[bbgemm.scala 846:22]
  assign st_27_io_GepAddr_valid = Gep_arrayidx2524_io_Out_1_valid; // @[bbgemm.scala 812:20]
  assign st_27_io_GepAddr_bits_data = Gep_arrayidx2524_io_Out_1_bits_data; // @[bbgemm.scala 812:20]
  assign st_27_io_inData_valid = FP_add2626_io_Out_0_valid; // @[bbgemm.scala 816:19]
  assign st_27_io_inData_bits_data = FP_add2626_io_Out_0_bits_data; // @[bbgemm.scala 816:19]
  assign st_27_io_MemReq_ready = MemCtrl_io_wr_mem_0_MemReq_ready; // @[bbgemm.scala 719:31]
  assign st_27_io_MemResp_valid = MemCtrl_io_wr_mem_0_MemResp_valid; // @[bbgemm.scala 721:20]
  assign binaryOp_indvars_iv_next28_clock = clock;
  assign binaryOp_indvars_iv_next28_reset = reset;
  assign binaryOp_indvars_iv_next28_io_enable_valid = bb_for_body165_io_Out_15_valid; // @[bbgemm.scala 615:40]
  assign binaryOp_indvars_iv_next28_io_enable_bits_taskID = bb_for_body165_io_Out_15_bits_taskID; // @[bbgemm.scala 615:40]
  assign binaryOp_indvars_iv_next28_io_enable_bits_control = bb_for_body165_io_Out_15_bits_control; // @[bbgemm.scala 615:40]
  assign binaryOp_indvars_iv_next28_io_Out_0_ready = Loop_0_io_CarryDepenIn_0_ready; // @[bbgemm.scala 481:29]
  assign binaryOp_indvars_iv_next28_io_Out_1_ready = icmp_exitcond29_io_LeftIO_ready; // @[bbgemm.scala 818:29]
  assign binaryOp_indvars_iv_next28_io_LeftIO_valid = phiindvars_iv16_io_Out_2_valid; // @[bbgemm.scala 794:40]
  assign binaryOp_indvars_iv_next28_io_LeftIO_bits_data = phiindvars_iv16_io_Out_2_bits_data; // @[bbgemm.scala 794:40]
  assign binaryOp_indvars_iv_next28_io_RightIO_valid = const7_io_Out_valid; // @[bbgemm.scala 748:41]
  assign icmp_exitcond29_clock = clock;
  assign icmp_exitcond29_reset = reset;
  assign icmp_exitcond29_io_enable_valid = bb_for_body165_io_Out_16_valid; // @[bbgemm.scala 618:29]
  assign icmp_exitcond29_io_enable_bits_taskID = bb_for_body165_io_Out_16_bits_taskID; // @[bbgemm.scala 618:29]
  assign icmp_exitcond29_io_enable_bits_control = bb_for_body165_io_Out_16_bits_control; // @[bbgemm.scala 618:29]
  assign icmp_exitcond29_io_Out_0_ready = br_30_io_CmpIO_ready; // @[bbgemm.scala 820:18]
  assign icmp_exitcond29_io_LeftIO_valid = binaryOp_indvars_iv_next28_io_Out_1_valid; // @[bbgemm.scala 818:29]
  assign icmp_exitcond29_io_LeftIO_bits_data = binaryOp_indvars_iv_next28_io_Out_1_bits_data; // @[bbgemm.scala 818:29]
  assign icmp_exitcond29_io_RightIO_valid = const8_io_Out_valid; // @[bbgemm.scala 750:30]
  assign br_30_clock = clock;
  assign br_30_reset = reset;
  assign br_30_io_enable_valid = bb_for_body165_io_Out_17_valid; // @[bbgemm.scala 621:19]
  assign br_30_io_enable_bits_taskID = bb_for_body165_io_Out_17_bits_taskID; // @[bbgemm.scala 621:19]
  assign br_30_io_enable_bits_control = bb_for_body165_io_Out_17_bits_control; // @[bbgemm.scala 621:19]
  assign br_30_io_CmpIO_valid = icmp_exitcond29_io_Out_0_valid; // @[bbgemm.scala 820:18]
  assign br_30_io_CmpIO_bits_taskID = icmp_exitcond29_io_Out_0_bits_taskID; // @[bbgemm.scala 820:18]
  assign br_30_io_CmpIO_bits_data = icmp_exitcond29_io_Out_0_bits_data; // @[bbgemm.scala 820:18]
  assign br_30_io_PredOp_0_valid = st_27_io_SuccOp_0_valid; // @[bbgemm.scala 846:22]
  assign br_30_io_TrueOutput_0_ready = Loop_0_io_loopFinish_0_ready; // @[bbgemm.scala 349:27]
  assign br_30_io_FalseOutput_0_ready = Loop_0_io_loopBack_0_ready; // @[bbgemm.scala 347:25]
  assign binaryOp_indvars_iv_next7231_clock = clock;
  assign binaryOp_indvars_iv_next7231_reset = reset;
  assign binaryOp_indvars_iv_next7231_io_enable_valid = bb_for_inc276_io_Out_2_valid; // @[bbgemm.scala 628:42]
  assign binaryOp_indvars_iv_next7231_io_enable_bits_taskID = bb_for_inc276_io_Out_2_bits_taskID; // @[bbgemm.scala 628:42]
  assign binaryOp_indvars_iv_next7231_io_enable_bits_control = bb_for_inc276_io_Out_2_bits_control; // @[bbgemm.scala 628:42]
  assign binaryOp_indvars_iv_next7231_io_Out_0_ready = Loop_1_io_CarryDepenIn_0_ready; // @[bbgemm.scala 483:29]
  assign binaryOp_indvars_iv_next7231_io_Out_1_ready = icmp_exitcond7732_io_LeftIO_ready; // @[bbgemm.scala 822:31]
  assign binaryOp_indvars_iv_next7231_io_LeftIO_valid = phiindvars_iv718_io_Out_2_valid; // @[bbgemm.scala 780:42]
  assign binaryOp_indvars_iv_next7231_io_LeftIO_bits_data = phiindvars_iv718_io_Out_2_bits_data; // @[bbgemm.scala 780:42]
  assign binaryOp_indvars_iv_next7231_io_RightIO_valid = const9_io_Out_valid; // @[bbgemm.scala 752:43]
  assign icmp_exitcond7732_clock = clock;
  assign icmp_exitcond7732_reset = reset;
  assign icmp_exitcond7732_io_enable_valid = bb_for_inc276_io_Out_3_valid; // @[bbgemm.scala 631:31]
  assign icmp_exitcond7732_io_enable_bits_taskID = bb_for_inc276_io_Out_3_bits_taskID; // @[bbgemm.scala 631:31]
  assign icmp_exitcond7732_io_enable_bits_control = bb_for_inc276_io_Out_3_bits_control; // @[bbgemm.scala 631:31]
  assign icmp_exitcond7732_io_Out_0_ready = br_33_io_CmpIO_ready; // @[bbgemm.scala 824:18]
  assign icmp_exitcond7732_io_LeftIO_valid = binaryOp_indvars_iv_next7231_io_Out_1_valid; // @[bbgemm.scala 822:31]
  assign icmp_exitcond7732_io_LeftIO_bits_data = binaryOp_indvars_iv_next7231_io_Out_1_bits_data; // @[bbgemm.scala 822:31]
  assign icmp_exitcond7732_io_RightIO_valid = const10_io_Out_valid; // @[bbgemm.scala 754:32]
  assign br_33_clock = clock;
  assign br_33_reset = reset;
  assign br_33_io_enable_valid = bb_for_inc276_io_Out_4_valid; // @[bbgemm.scala 634:19]
  assign br_33_io_enable_bits_taskID = bb_for_inc276_io_Out_4_bits_taskID; // @[bbgemm.scala 634:19]
  assign br_33_io_enable_bits_control = bb_for_inc276_io_Out_4_bits_control; // @[bbgemm.scala 634:19]
  assign br_33_io_CmpIO_valid = icmp_exitcond7732_io_Out_0_valid; // @[bbgemm.scala 824:18]
  assign br_33_io_CmpIO_bits_taskID = icmp_exitcond7732_io_Out_0_bits_taskID; // @[bbgemm.scala 824:18]
  assign br_33_io_CmpIO_bits_data = icmp_exitcond7732_io_Out_0_bits_data; // @[bbgemm.scala 824:18]
  assign br_33_io_TrueOutput_0_ready = Loop_1_io_loopFinish_0_ready; // @[bbgemm.scala 355:27]
  assign br_33_io_FalseOutput_0_ready = Loop_1_io_loopBack_0_ready; // @[bbgemm.scala 353:25]
  assign binaryOp_indvars_iv_next7934_clock = clock;
  assign binaryOp_indvars_iv_next7934_reset = reset;
  assign binaryOp_indvars_iv_next7934_io_enable_valid = bb_for_inc307_io_Out_2_valid; // @[bbgemm.scala 641:42]
  assign binaryOp_indvars_iv_next7934_io_enable_bits_taskID = bb_for_inc307_io_Out_2_bits_taskID; // @[bbgemm.scala 641:42]
  assign binaryOp_indvars_iv_next7934_io_enable_bits_control = bb_for_inc307_io_Out_2_bits_control; // @[bbgemm.scala 641:42]
  assign binaryOp_indvars_iv_next7934_io_Out_0_ready = Loop_2_io_CarryDepenIn_0_ready; // @[bbgemm.scala 485:29]
  assign binaryOp_indvars_iv_next7934_io_Out_1_ready = icmp_exitcond8135_io_LeftIO_ready; // @[bbgemm.scala 826:31]
  assign binaryOp_indvars_iv_next7934_io_LeftIO_valid = phiindvars_iv785_io_Out_1_valid; // @[bbgemm.scala 774:42]
  assign binaryOp_indvars_iv_next7934_io_LeftIO_bits_data = phiindvars_iv785_io_Out_1_bits_data; // @[bbgemm.scala 774:42]
  assign binaryOp_indvars_iv_next7934_io_RightIO_valid = const11_io_Out_valid; // @[bbgemm.scala 756:43]
  assign icmp_exitcond8135_clock = clock;
  assign icmp_exitcond8135_reset = reset;
  assign icmp_exitcond8135_io_enable_valid = bb_for_inc307_io_Out_3_valid; // @[bbgemm.scala 644:31]
  assign icmp_exitcond8135_io_enable_bits_taskID = bb_for_inc307_io_Out_3_bits_taskID; // @[bbgemm.scala 644:31]
  assign icmp_exitcond8135_io_enable_bits_control = bb_for_inc307_io_Out_3_bits_control; // @[bbgemm.scala 644:31]
  assign icmp_exitcond8135_io_Out_0_ready = br_36_io_CmpIO_ready; // @[bbgemm.scala 828:18]
  assign icmp_exitcond8135_io_LeftIO_valid = binaryOp_indvars_iv_next7934_io_Out_1_valid; // @[bbgemm.scala 826:31]
  assign icmp_exitcond8135_io_LeftIO_bits_data = binaryOp_indvars_iv_next7934_io_Out_1_bits_data; // @[bbgemm.scala 826:31]
  assign icmp_exitcond8135_io_RightIO_valid = const12_io_Out_valid; // @[bbgemm.scala 758:32]
  assign br_36_clock = clock;
  assign br_36_reset = reset;
  assign br_36_io_enable_valid = bb_for_inc307_io_Out_4_valid; // @[bbgemm.scala 647:19]
  assign br_36_io_enable_bits_taskID = bb_for_inc307_io_Out_4_bits_taskID; // @[bbgemm.scala 647:19]
  assign br_36_io_enable_bits_control = bb_for_inc307_io_Out_4_bits_control; // @[bbgemm.scala 647:19]
  assign br_36_io_CmpIO_valid = icmp_exitcond8135_io_Out_0_valid; // @[bbgemm.scala 828:18]
  assign br_36_io_CmpIO_bits_taskID = icmp_exitcond8135_io_Out_0_bits_taskID; // @[bbgemm.scala 828:18]
  assign br_36_io_CmpIO_bits_data = icmp_exitcond8135_io_Out_0_bits_data; // @[bbgemm.scala 828:18]
  assign br_36_io_TrueOutput_0_ready = Loop_2_io_loopFinish_0_ready; // @[bbgemm.scala 361:27]
  assign br_36_io_FalseOutput_0_ready = Loop_2_io_loopBack_0_ready; // @[bbgemm.scala 359:25]
  assign binaryOp_indvars_iv_next8337_clock = clock;
  assign binaryOp_indvars_iv_next8337_reset = reset;
  assign binaryOp_indvars_iv_next8337_io_enable_valid = bb_for_inc338_io_Out_2_valid; // @[bbgemm.scala 654:42]
  assign binaryOp_indvars_iv_next8337_io_enable_bits_taskID = bb_for_inc338_io_Out_2_bits_taskID; // @[bbgemm.scala 654:42]
  assign binaryOp_indvars_iv_next8337_io_enable_bits_control = bb_for_inc338_io_Out_2_bits_control; // @[bbgemm.scala 654:42]
  assign binaryOp_indvars_iv_next8337_io_Out_0_ready = Loop_3_io_CarryDepenIn_0_ready; // @[bbgemm.scala 487:29]
  assign binaryOp_indvars_iv_next8337_io_Out_1_ready = icmp_cmp238_io_LeftIO_ready; // @[bbgemm.scala 830:25]
  assign binaryOp_indvars_iv_next8337_io_LeftIO_valid = phiindvars_iv823_io_Out_1_valid; // @[bbgemm.scala 770:42]
  assign binaryOp_indvars_iv_next8337_io_LeftIO_bits_data = phiindvars_iv823_io_Out_1_bits_data; // @[bbgemm.scala 770:42]
  assign binaryOp_indvars_iv_next8337_io_RightIO_valid = const13_io_Out_valid; // @[bbgemm.scala 760:43]
  assign icmp_cmp238_clock = clock;
  assign icmp_cmp238_reset = reset;
  assign icmp_cmp238_io_enable_valid = bb_for_inc338_io_Out_3_valid; // @[bbgemm.scala 657:25]
  assign icmp_cmp238_io_enable_bits_taskID = bb_for_inc338_io_Out_3_bits_taskID; // @[bbgemm.scala 657:25]
  assign icmp_cmp238_io_enable_bits_control = bb_for_inc338_io_Out_3_bits_control; // @[bbgemm.scala 657:25]
  assign icmp_cmp238_io_Out_0_ready = br_39_io_CmpIO_ready; // @[bbgemm.scala 832:18]
  assign icmp_cmp238_io_LeftIO_valid = binaryOp_indvars_iv_next8337_io_Out_1_valid; // @[bbgemm.scala 830:25]
  assign icmp_cmp238_io_LeftIO_bits_data = binaryOp_indvars_iv_next8337_io_Out_1_bits_data; // @[bbgemm.scala 830:25]
  assign icmp_cmp238_io_RightIO_valid = const14_io_Out_valid; // @[bbgemm.scala 762:26]
  assign br_39_clock = clock;
  assign br_39_reset = reset;
  assign br_39_io_enable_valid = bb_for_inc338_io_Out_4_valid; // @[bbgemm.scala 660:19]
  assign br_39_io_enable_bits_taskID = bb_for_inc338_io_Out_4_bits_taskID; // @[bbgemm.scala 660:19]
  assign br_39_io_enable_bits_control = bb_for_inc338_io_Out_4_bits_control; // @[bbgemm.scala 660:19]
  assign br_39_io_CmpIO_valid = icmp_cmp238_io_Out_0_valid; // @[bbgemm.scala 832:18]
  assign br_39_io_CmpIO_bits_taskID = icmp_cmp238_io_Out_0_bits_taskID; // @[bbgemm.scala 832:18]
  assign br_39_io_CmpIO_bits_data = icmp_cmp238_io_Out_0_bits_data; // @[bbgemm.scala 832:18]
  assign br_39_io_TrueOutput_0_ready = Loop_3_io_loopBack_0_ready; // @[bbgemm.scala 365:25]
  assign br_39_io_FalseOutput_0_ready = Loop_3_io_loopFinish_0_ready; // @[bbgemm.scala 367:27]
  assign binaryOp_indvars_iv_next8540_clock = clock;
  assign binaryOp_indvars_iv_next8540_reset = reset;
  assign binaryOp_indvars_iv_next8540_io_enable_valid = bb_for_inc369_io_Out_2_valid; // @[bbgemm.scala 667:42]
  assign binaryOp_indvars_iv_next8540_io_enable_bits_taskID = bb_for_inc369_io_Out_2_bits_taskID; // @[bbgemm.scala 667:42]
  assign binaryOp_indvars_iv_next8540_io_enable_bits_control = bb_for_inc369_io_Out_2_bits_control; // @[bbgemm.scala 667:42]
  assign binaryOp_indvars_iv_next8540_io_Out_0_ready = Loop_4_io_CarryDepenIn_0_ready; // @[bbgemm.scala 489:29]
  assign binaryOp_indvars_iv_next8540_io_Out_1_ready = icmp_cmp41_io_LeftIO_ready; // @[bbgemm.scala 834:24]
  assign binaryOp_indvars_iv_next8540_io_LeftIO_valid = phiindvars_iv841_io_Out_1_valid; // @[bbgemm.scala 768:42]
  assign binaryOp_indvars_iv_next8540_io_LeftIO_bits_data = phiindvars_iv841_io_Out_1_bits_data; // @[bbgemm.scala 768:42]
  assign binaryOp_indvars_iv_next8540_io_RightIO_valid = const15_io_Out_valid; // @[bbgemm.scala 764:43]
  assign icmp_cmp41_clock = clock;
  assign icmp_cmp41_reset = reset;
  assign icmp_cmp41_io_enable_valid = bb_for_inc369_io_Out_3_valid; // @[bbgemm.scala 670:24]
  assign icmp_cmp41_io_enable_bits_taskID = bb_for_inc369_io_Out_3_bits_taskID; // @[bbgemm.scala 670:24]
  assign icmp_cmp41_io_enable_bits_control = bb_for_inc369_io_Out_3_bits_control; // @[bbgemm.scala 670:24]
  assign icmp_cmp41_io_Out_0_ready = br_42_io_CmpIO_ready; // @[bbgemm.scala 836:18]
  assign icmp_cmp41_io_LeftIO_valid = binaryOp_indvars_iv_next8540_io_Out_1_valid; // @[bbgemm.scala 834:24]
  assign icmp_cmp41_io_LeftIO_bits_data = binaryOp_indvars_iv_next8540_io_Out_1_bits_data; // @[bbgemm.scala 834:24]
  assign icmp_cmp41_io_RightIO_valid = const16_io_Out_valid; // @[bbgemm.scala 766:25]
  assign br_42_clock = clock;
  assign br_42_reset = reset;
  assign br_42_io_enable_valid = bb_for_inc369_io_Out_4_valid; // @[bbgemm.scala 673:19]
  assign br_42_io_enable_bits_taskID = bb_for_inc369_io_Out_4_bits_taskID; // @[bbgemm.scala 673:19]
  assign br_42_io_enable_bits_control = bb_for_inc369_io_Out_4_bits_control; // @[bbgemm.scala 673:19]
  assign br_42_io_CmpIO_valid = icmp_cmp41_io_Out_0_valid; // @[bbgemm.scala 836:18]
  assign br_42_io_CmpIO_bits_taskID = icmp_cmp41_io_Out_0_bits_taskID; // @[bbgemm.scala 836:18]
  assign br_42_io_CmpIO_bits_data = icmp_cmp41_io_Out_0_bits_data; // @[bbgemm.scala 836:18]
  assign br_42_io_TrueOutput_0_ready = Loop_4_io_loopBack_0_ready; // @[bbgemm.scala 371:25]
  assign br_42_io_FalseOutput_0_ready = Loop_4_io_loopFinish_0_ready; // @[bbgemm.scala 373:27]
  assign ret_43_clock = clock;
  assign ret_43_reset = reset;
  assign ret_43_io_In_enable_valid = bb_for_end3810_io_Out_0_valid; // @[bbgemm.scala 676:23]
  assign ret_43_io_In_enable_bits_taskID = bb_for_end3810_io_Out_0_bits_taskID; // @[bbgemm.scala 676:23]
  assign ret_43_io_Out_ready = io_out_ready; // @[bbgemm.scala 854:10]
  assign const0_clock = clock;
  assign const0_reset = reset;
  assign const0_io_enable_valid = bb_loopkk1_io_Out_0_valid; // @[bbgemm.scala 516:20]
  assign const0_io_enable_bits_taskID = bb_loopkk1_io_Out_0_bits_taskID; // @[bbgemm.scala 516:20]
  assign const0_io_enable_bits_control = bb_loopkk1_io_Out_0_bits_control; // @[bbgemm.scala 516:20]
  assign const0_io_Out_ready = phiindvars_iv841_io_InData_0_ready; // @[bbgemm.scala 734:33]
  assign const1_clock = clock;
  assign const1_reset = reset;
  assign const1_io_enable_valid = bb_loopi2_io_Out_0_valid; // @[bbgemm.scala 524:20]
  assign const1_io_enable_bits_taskID = bb_loopi2_io_Out_0_bits_taskID; // @[bbgemm.scala 524:20]
  assign const1_io_enable_bits_control = bb_loopi2_io_Out_0_bits_control; // @[bbgemm.scala 524:20]
  assign const1_io_Out_ready = phiindvars_iv823_io_InData_0_ready; // @[bbgemm.scala 736:33]
  assign const2_clock = clock;
  assign const2_reset = reset;
  assign const2_io_enable_valid = bb_loopk3_io_Out_0_valid; // @[bbgemm.scala 532:20]
  assign const2_io_enable_bits_taskID = bb_loopk3_io_Out_0_bits_taskID; // @[bbgemm.scala 532:20]
  assign const2_io_enable_bits_control = bb_loopk3_io_Out_0_bits_control; // @[bbgemm.scala 532:20]
  assign const2_io_Out_ready = phiindvars_iv785_io_InData_0_ready; // @[bbgemm.scala 738:33]
  assign const3_clock = clock;
  assign const3_reset = reset;
  assign const3_io_enable_valid = bb_loopk3_io_Out_1_valid; // @[bbgemm.scala 534:20]
  assign const3_io_enable_bits_taskID = bb_loopk3_io_Out_1_bits_taskID; // @[bbgemm.scala 534:20]
  assign const3_io_enable_bits_control = bb_loopk3_io_Out_1_bits_control; // @[bbgemm.scala 534:20]
  assign const3_io_Out_ready = binaryOp_6_io_RightIO_ready; // @[bbgemm.scala 740:25]
  assign const4_clock = clock;
  assign const4_reset = reset;
  assign const4_io_enable_valid = bb_for_body94_io_Out_0_valid; // @[bbgemm.scala 545:20]
  assign const4_io_enable_bits_taskID = bb_for_body94_io_Out_0_bits_taskID; // @[bbgemm.scala 545:20]
  assign const4_io_enable_bits_control = bb_for_body94_io_Out_0_bits_control; // @[bbgemm.scala 545:20]
  assign const4_io_Out_ready = phiindvars_iv718_io_InData_0_ready; // @[bbgemm.scala 742:33]
  assign const5_clock = clock;
  assign const5_reset = reset;
  assign const5_io_enable_valid = bb_for_body94_io_Out_1_valid; // @[bbgemm.scala 547:20]
  assign const5_io_enable_bits_taskID = bb_for_body94_io_Out_1_bits_taskID; // @[bbgemm.scala 547:20]
  assign const5_io_enable_bits_control = bb_for_body94_io_Out_1_bits_control; // @[bbgemm.scala 547:20]
  assign const5_io_Out_ready = binaryOp_10_io_RightIO_ready; // @[bbgemm.scala 744:26]
  assign const6_clock = clock;
  assign const6_reset = reset;
  assign const6_io_enable_valid = bb_for_body165_io_Out_0_valid; // @[bbgemm.scala 573:20]
  assign const6_io_enable_bits_taskID = bb_for_body165_io_Out_0_bits_taskID; // @[bbgemm.scala 573:20]
  assign const6_io_enable_bits_control = bb_for_body165_io_Out_0_bits_control; // @[bbgemm.scala 573:20]
  assign const6_io_Out_ready = phiindvars_iv16_io_InData_0_ready; // @[bbgemm.scala 746:32]
  assign const7_clock = clock;
  assign const7_reset = reset;
  assign const7_io_enable_valid = bb_for_body165_io_Out_1_valid; // @[bbgemm.scala 575:20]
  assign const7_io_enable_bits_taskID = bb_for_body165_io_Out_1_bits_taskID; // @[bbgemm.scala 575:20]
  assign const7_io_enable_bits_control = bb_for_body165_io_Out_1_bits_control; // @[bbgemm.scala 575:20]
  assign const7_io_Out_ready = binaryOp_indvars_iv_next28_io_RightIO_ready; // @[bbgemm.scala 748:41]
  assign const8_clock = clock;
  assign const8_reset = reset;
  assign const8_io_enable_valid = bb_for_body165_io_Out_2_valid; // @[bbgemm.scala 577:20]
  assign const8_io_enable_bits_taskID = bb_for_body165_io_Out_2_bits_taskID; // @[bbgemm.scala 577:20]
  assign const8_io_enable_bits_control = bb_for_body165_io_Out_2_bits_control; // @[bbgemm.scala 577:20]
  assign const8_io_Out_ready = icmp_exitcond29_io_RightIO_ready; // @[bbgemm.scala 750:30]
  assign const9_clock = clock;
  assign const9_reset = reset;
  assign const9_io_enable_valid = bb_for_inc276_io_Out_0_valid; // @[bbgemm.scala 624:20]
  assign const9_io_enable_bits_taskID = bb_for_inc276_io_Out_0_bits_taskID; // @[bbgemm.scala 624:20]
  assign const9_io_enable_bits_control = bb_for_inc276_io_Out_0_bits_control; // @[bbgemm.scala 624:20]
  assign const9_io_Out_ready = binaryOp_indvars_iv_next7231_io_RightIO_ready; // @[bbgemm.scala 752:43]
  assign const10_clock = clock;
  assign const10_reset = reset;
  assign const10_io_enable_valid = bb_for_inc276_io_Out_1_valid; // @[bbgemm.scala 626:21]
  assign const10_io_enable_bits_taskID = bb_for_inc276_io_Out_1_bits_taskID; // @[bbgemm.scala 626:21]
  assign const10_io_enable_bits_control = bb_for_inc276_io_Out_1_bits_control; // @[bbgemm.scala 626:21]
  assign const10_io_Out_ready = icmp_exitcond7732_io_RightIO_ready; // @[bbgemm.scala 754:32]
  assign const11_clock = clock;
  assign const11_reset = reset;
  assign const11_io_enable_valid = bb_for_inc307_io_Out_0_valid; // @[bbgemm.scala 637:21]
  assign const11_io_enable_bits_taskID = bb_for_inc307_io_Out_0_bits_taskID; // @[bbgemm.scala 637:21]
  assign const11_io_enable_bits_control = bb_for_inc307_io_Out_0_bits_control; // @[bbgemm.scala 637:21]
  assign const11_io_Out_ready = binaryOp_indvars_iv_next7934_io_RightIO_ready; // @[bbgemm.scala 756:43]
  assign const12_clock = clock;
  assign const12_reset = reset;
  assign const12_io_enable_valid = bb_for_inc307_io_Out_1_valid; // @[bbgemm.scala 639:21]
  assign const12_io_enable_bits_taskID = bb_for_inc307_io_Out_1_bits_taskID; // @[bbgemm.scala 639:21]
  assign const12_io_enable_bits_control = bb_for_inc307_io_Out_1_bits_control; // @[bbgemm.scala 639:21]
  assign const12_io_Out_ready = icmp_exitcond8135_io_RightIO_ready; // @[bbgemm.scala 758:32]
  assign const13_clock = clock;
  assign const13_reset = reset;
  assign const13_io_enable_valid = bb_for_inc338_io_Out_0_valid; // @[bbgemm.scala 650:21]
  assign const13_io_enable_bits_taskID = bb_for_inc338_io_Out_0_bits_taskID; // @[bbgemm.scala 650:21]
  assign const13_io_enable_bits_control = bb_for_inc338_io_Out_0_bits_control; // @[bbgemm.scala 650:21]
  assign const13_io_Out_ready = binaryOp_indvars_iv_next8337_io_RightIO_ready; // @[bbgemm.scala 760:43]
  assign const14_clock = clock;
  assign const14_reset = reset;
  assign const14_io_enable_valid = bb_for_inc338_io_Out_1_valid; // @[bbgemm.scala 652:21]
  assign const14_io_enable_bits_taskID = bb_for_inc338_io_Out_1_bits_taskID; // @[bbgemm.scala 652:21]
  assign const14_io_enable_bits_control = bb_for_inc338_io_Out_1_bits_control; // @[bbgemm.scala 652:21]
  assign const14_io_Out_ready = icmp_cmp238_io_RightIO_ready; // @[bbgemm.scala 762:26]
  assign const15_clock = clock;
  assign const15_reset = reset;
  assign const15_io_enable_valid = bb_for_inc369_io_Out_0_valid; // @[bbgemm.scala 663:21]
  assign const15_io_enable_bits_taskID = bb_for_inc369_io_Out_0_bits_taskID; // @[bbgemm.scala 663:21]
  assign const15_io_enable_bits_control = bb_for_inc369_io_Out_0_bits_control; // @[bbgemm.scala 663:21]
  assign const15_io_Out_ready = binaryOp_indvars_iv_next8540_io_RightIO_ready; // @[bbgemm.scala 764:43]
  assign const16_clock = clock;
  assign const16_reset = reset;
  assign const16_io_enable_valid = bb_for_inc369_io_Out_1_valid; // @[bbgemm.scala 665:21]
  assign const16_io_enable_bits_taskID = bb_for_inc369_io_Out_1_bits_taskID; // @[bbgemm.scala 665:21]
  assign const16_io_enable_bits_control = bb_for_inc369_io_Out_1_bits_control; // @[bbgemm.scala 665:21]
  assign const16_io_Out_ready = icmp_cmp41_io_RightIO_ready; // @[bbgemm.scala 766:25]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  input         io_enq_valid,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits,
  output [1:0]  io_count
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram [0:1]; // @[Decoupled.scala 218:16]
  wire [63:0] ram__T_11_data; // @[Decoupled.scala 218:16]
  wire  ram__T_11_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram__T_3_data; // @[Decoupled.scala 218:16]
  wire  ram__T_3_addr; // @[Decoupled.scala 218:16]
  wire  ram__T_3_mask; // @[Decoupled.scala 218:16]
  wire  ram__T_3_en; // @[Decoupled.scala 218:16]
  reg  deq_ptr_value; // @[Counter.scala 29:33]
  wire  ptr_match = ~deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = deq_ptr_value + 1'h1; // @[Counter.scala 39:22]
  wire  ptr_diff = 1'h0 - deq_ptr_value; // @[Decoupled.scala 257:32]
  assign ram__T_11_addr = deq_ptr_value;
  assign ram__T_11_data = ram[ram__T_11_addr]; // @[Decoupled.scala 218:16]
  assign ram__T_3_data = 64'h0;
  assign ram__T_3_addr = 1'h0;
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = 1'h0;
  assign io_deq_valid = ~ptr_match; // @[Decoupled.scala 240:16]
  assign io_deq_bits = ram__T_11_data; // @[Decoupled.scala 242:15]
  assign io_count = {{1'd0}, ptr_diff}; // @[Decoupled.scala 259:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  deq_ptr_value = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin
      deq_ptr_value <= 1'h0;
    end else if (do_deq) begin
      deq_ptr_value <= _T_7;
    end
  end
endmodule
module DebugVMEBufferNode(
  input         clock,
  input         reset,
  input  [31:0] io_addrDebug,
  input         io_vmeOut_cmd_ready,
  output        io_vmeOut_cmd_valid,
  output [31:0] io_vmeOut_cmd_bits_addr,
  output [7:0]  io_vmeOut_cmd_bits_len,
  input         io_vmeOut_data_ready,
  output        io_vmeOut_data_valid,
  output [63:0] io_vmeOut_data_bits,
  input         io_vmeOut_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  LogData_clock; // @[DebugStore.scala 243:23]
  wire  LogData_reset; // @[DebugStore.scala 243:23]
  wire  LogData_io_enq_valid; // @[DebugStore.scala 243:23]
  wire  LogData_io_deq_ready; // @[DebugStore.scala 243:23]
  wire  LogData_io_deq_valid; // @[DebugStore.scala 243:23]
  wire [63:0] LogData_io_deq_bits; // @[DebugStore.scala 243:23]
  wire [1:0] LogData_io_count; // @[DebugStore.scala 243:23]
  reg [63:0] addr_debug_reg; // @[DebugStore.scala 238:31]
  reg [1:0] wState; // @[DebugStore.scala 240:23]
  reg  queue_count; // @[DebugStore.scala 246:28]
  wire  _T_4 = LogData_io_enq_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = queue_count + 1'h1; // @[DebugStore.scala 248:32]
  wire [63:0] _GEN_20 = {{32'd0}, io_addrDebug}; // @[DebugStore.scala 259:43]
  wire [63:0] _T_13 = _GEN_20 + addr_debug_reg; // @[DebugStore.scala 259:43]
  wire  _T_15 = queue_count - 1'h1; // @[DebugStore.scala 260:41]
  wire  _T_17 = 2'h0 == wState; // @[Conditional.scala 37:30]
  wire  _T_20 = LogData_io_count == 2'h1; // @[DebugStore.scala 266:82]
  wire  _T_22 = 2'h1 == wState; // @[Conditional.scala 37:30]
  wire  _T_23 = io_vmeOut_cmd_ready & io_vmeOut_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _T_24 = 2'h2 == wState; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_21 = {{3'd0}, queue_count}; // @[DebugStore.scala 279:57]
  wire [4:0] _T_25 = _GEN_21 * 4'h8; // @[DebugStore.scala 279:57]
  wire [63:0] _GEN_22 = {{59'd0}, _T_25}; // @[DebugStore.scala 279:42]
  wire [63:0] _T_27 = addr_debug_reg + _GEN_22; // @[DebugStore.scala 279:42]
  wire  _T_28 = wState == 2'h2; // @[DebugStore.scala 289:15]
  Queue_3 LogData ( // @[DebugStore.scala 243:23]
    .clock(LogData_clock),
    .reset(LogData_reset),
    .io_enq_valid(LogData_io_enq_valid),
    .io_deq_ready(LogData_io_deq_ready),
    .io_deq_valid(LogData_io_deq_valid),
    .io_deq_bits(LogData_io_deq_bits),
    .io_count(LogData_io_count)
  );
  assign io_vmeOut_cmd_valid = wState == 2'h1; // @[DebugStore.scala 261:23]
  assign io_vmeOut_cmd_bits_addr = _T_13[31:0]; // @[DebugStore.scala 259:27]
  assign io_vmeOut_cmd_bits_len = {{7'd0}, _T_15}; // @[DebugStore.scala 260:26]
  assign io_vmeOut_data_valid = _T_28 & LogData_io_deq_valid; // @[DebugStore.scala 286:24 DebugStore.scala 291:26]
  assign io_vmeOut_data_bits = _T_28 ? LogData_io_deq_bits : 64'h0; // @[DebugStore.scala 285:23 DebugStore.scala 290:25]
  assign LogData_clock = clock;
  assign LogData_reset = reset;
  assign LogData_io_enq_valid = 1'h0; // @[DebugStore.scala 256:24]
  assign LogData_io_deq_ready = _T_28 & io_vmeOut_data_ready; // @[DebugStore.scala 287:24 DebugStore.scala 292:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addr_debug_reg = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  wState = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  queue_count = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      addr_debug_reg <= 64'h0;
    end else if (!(_T_17)) begin
      if (!(_T_22)) begin
        if (_T_24) begin
          if (io_vmeOut_ack) begin
            addr_debug_reg <= _T_27;
          end
        end
      end
    end
    if (reset) begin
      wState <= 2'h0;
    end else if (_T_17) begin
      if (_T_20) begin
        wState <= 2'h1;
      end
    end else if (_T_22) begin
      if (_T_23) begin
        wState <= 2'h2;
      end
    end else if (_T_24) begin
      if (io_vmeOut_ack) begin
        wState <= 2'h0;
      end
    end
    if (reset) begin
      queue_count <= 1'h0;
    end else if (_T_17) begin
      if (_T_4) begin
        queue_count <= _T_6;
      end
    end else if (_T_22) begin
      if (_T_4) begin
        queue_count <= _T_6;
      end
    end else if (_T_24) begin
      if (io_vmeOut_ack) begin
        queue_count <= 1'h0;
      end else if (_T_4) begin
        queue_count <= _T_6;
      end
    end else if (_T_4) begin
      queue_count <= _T_6;
    end
  end
endmodule
module DebugBufferWriters(
  input         clock,
  input         reset,
  input  [31:0] io_addrDebug_0,
  input  [31:0] io_addrDebug_1,
  input  [31:0] io_addrDebug_2,
  input         io_vmeOut_0_cmd_ready,
  output        io_vmeOut_0_cmd_valid,
  output [31:0] io_vmeOut_0_cmd_bits_addr,
  output [7:0]  io_vmeOut_0_cmd_bits_len,
  input         io_vmeOut_0_data_ready,
  output        io_vmeOut_0_data_valid,
  output [63:0] io_vmeOut_0_data_bits,
  input         io_vmeOut_0_ack,
  input         io_vmeOut_1_cmd_ready,
  output        io_vmeOut_1_cmd_valid,
  output [31:0] io_vmeOut_1_cmd_bits_addr,
  output [7:0]  io_vmeOut_1_cmd_bits_len,
  input         io_vmeOut_1_data_ready,
  output        io_vmeOut_1_data_valid,
  output [63:0] io_vmeOut_1_data_bits,
  input         io_vmeOut_1_ack,
  input         io_vmeOut_2_cmd_ready,
  output        io_vmeOut_2_cmd_valid,
  output [31:0] io_vmeOut_2_cmd_bits_addr,
  output [7:0]  io_vmeOut_2_cmd_bits_len,
  input         io_vmeOut_2_data_ready,
  output        io_vmeOut_2_data_valid,
  output [63:0] io_vmeOut_2_data_bits,
  input         io_vmeOut_2_ack
);
  wire  buffers_0_clock; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_0_reset; // @[DebugBufferWriters.scala 23:52]
  wire [31:0] buffers_0_io_addrDebug; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_0_io_vmeOut_cmd_ready; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_0_io_vmeOut_cmd_valid; // @[DebugBufferWriters.scala 23:52]
  wire [31:0] buffers_0_io_vmeOut_cmd_bits_addr; // @[DebugBufferWriters.scala 23:52]
  wire [7:0] buffers_0_io_vmeOut_cmd_bits_len; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_0_io_vmeOut_data_ready; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_0_io_vmeOut_data_valid; // @[DebugBufferWriters.scala 23:52]
  wire [63:0] buffers_0_io_vmeOut_data_bits; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_0_io_vmeOut_ack; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_clock; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_reset; // @[DebugBufferWriters.scala 23:52]
  wire [31:0] buffers_1_io_addrDebug; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_io_vmeOut_cmd_ready; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_io_vmeOut_cmd_valid; // @[DebugBufferWriters.scala 23:52]
  wire [31:0] buffers_1_io_vmeOut_cmd_bits_addr; // @[DebugBufferWriters.scala 23:52]
  wire [7:0] buffers_1_io_vmeOut_cmd_bits_len; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_io_vmeOut_data_ready; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_io_vmeOut_data_valid; // @[DebugBufferWriters.scala 23:52]
  wire [63:0] buffers_1_io_vmeOut_data_bits; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_1_io_vmeOut_ack; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_clock; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_reset; // @[DebugBufferWriters.scala 23:52]
  wire [31:0] buffers_2_io_addrDebug; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_io_vmeOut_cmd_ready; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_io_vmeOut_cmd_valid; // @[DebugBufferWriters.scala 23:52]
  wire [31:0] buffers_2_io_vmeOut_cmd_bits_addr; // @[DebugBufferWriters.scala 23:52]
  wire [7:0] buffers_2_io_vmeOut_cmd_bits_len; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_io_vmeOut_data_ready; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_io_vmeOut_data_valid; // @[DebugBufferWriters.scala 23:52]
  wire [63:0] buffers_2_io_vmeOut_data_bits; // @[DebugBufferWriters.scala 23:52]
  wire  buffers_2_io_vmeOut_ack; // @[DebugBufferWriters.scala 23:52]
  DebugVMEBufferNode buffers_0 ( // @[DebugBufferWriters.scala 23:52]
    .clock(buffers_0_clock),
    .reset(buffers_0_reset),
    .io_addrDebug(buffers_0_io_addrDebug),
    .io_vmeOut_cmd_ready(buffers_0_io_vmeOut_cmd_ready),
    .io_vmeOut_cmd_valid(buffers_0_io_vmeOut_cmd_valid),
    .io_vmeOut_cmd_bits_addr(buffers_0_io_vmeOut_cmd_bits_addr),
    .io_vmeOut_cmd_bits_len(buffers_0_io_vmeOut_cmd_bits_len),
    .io_vmeOut_data_ready(buffers_0_io_vmeOut_data_ready),
    .io_vmeOut_data_valid(buffers_0_io_vmeOut_data_valid),
    .io_vmeOut_data_bits(buffers_0_io_vmeOut_data_bits),
    .io_vmeOut_ack(buffers_0_io_vmeOut_ack)
  );
  DebugVMEBufferNode buffers_1 ( // @[DebugBufferWriters.scala 23:52]
    .clock(buffers_1_clock),
    .reset(buffers_1_reset),
    .io_addrDebug(buffers_1_io_addrDebug),
    .io_vmeOut_cmd_ready(buffers_1_io_vmeOut_cmd_ready),
    .io_vmeOut_cmd_valid(buffers_1_io_vmeOut_cmd_valid),
    .io_vmeOut_cmd_bits_addr(buffers_1_io_vmeOut_cmd_bits_addr),
    .io_vmeOut_cmd_bits_len(buffers_1_io_vmeOut_cmd_bits_len),
    .io_vmeOut_data_ready(buffers_1_io_vmeOut_data_ready),
    .io_vmeOut_data_valid(buffers_1_io_vmeOut_data_valid),
    .io_vmeOut_data_bits(buffers_1_io_vmeOut_data_bits),
    .io_vmeOut_ack(buffers_1_io_vmeOut_ack)
  );
  DebugVMEBufferNode buffers_2 ( // @[DebugBufferWriters.scala 23:52]
    .clock(buffers_2_clock),
    .reset(buffers_2_reset),
    .io_addrDebug(buffers_2_io_addrDebug),
    .io_vmeOut_cmd_ready(buffers_2_io_vmeOut_cmd_ready),
    .io_vmeOut_cmd_valid(buffers_2_io_vmeOut_cmd_valid),
    .io_vmeOut_cmd_bits_addr(buffers_2_io_vmeOut_cmd_bits_addr),
    .io_vmeOut_cmd_bits_len(buffers_2_io_vmeOut_cmd_bits_len),
    .io_vmeOut_data_ready(buffers_2_io_vmeOut_data_ready),
    .io_vmeOut_data_valid(buffers_2_io_vmeOut_data_valid),
    .io_vmeOut_data_bits(buffers_2_io_vmeOut_data_bits),
    .io_vmeOut_ack(buffers_2_io_vmeOut_ack)
  );
  assign io_vmeOut_0_cmd_valid = buffers_0_io_vmeOut_cmd_valid; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_0_cmd_bits_addr = buffers_0_io_vmeOut_cmd_bits_addr; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_0_cmd_bits_len = buffers_0_io_vmeOut_cmd_bits_len; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_0_data_valid = buffers_0_io_vmeOut_data_valid; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_0_data_bits = buffers_0_io_vmeOut_data_bits; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_1_cmd_valid = buffers_1_io_vmeOut_cmd_valid; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_1_cmd_bits_addr = buffers_1_io_vmeOut_cmd_bits_addr; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_1_cmd_bits_len = buffers_1_io_vmeOut_cmd_bits_len; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_1_data_valid = buffers_1_io_vmeOut_data_valid; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_1_data_bits = buffers_1_io_vmeOut_data_bits; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_2_cmd_valid = buffers_2_io_vmeOut_cmd_valid; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_2_cmd_bits_addr = buffers_2_io_vmeOut_cmd_bits_addr; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_2_cmd_bits_len = buffers_2_io_vmeOut_cmd_bits_len; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_2_data_valid = buffers_2_io_vmeOut_data_valid; // @[DebugBufferWriters.scala 48:18]
  assign io_vmeOut_2_data_bits = buffers_2_io_vmeOut_data_bits; // @[DebugBufferWriters.scala 48:18]
  assign buffers_0_clock = clock;
  assign buffers_0_reset = reset;
  assign buffers_0_io_addrDebug = io_addrDebug_0; // @[DebugBufferWriters.scala 47:29]
  assign buffers_0_io_vmeOut_cmd_ready = io_vmeOut_0_cmd_ready; // @[DebugBufferWriters.scala 48:18]
  assign buffers_0_io_vmeOut_data_ready = io_vmeOut_0_data_ready; // @[DebugBufferWriters.scala 48:18]
  assign buffers_0_io_vmeOut_ack = io_vmeOut_0_ack; // @[DebugBufferWriters.scala 48:18]
  assign buffers_1_clock = clock;
  assign buffers_1_reset = reset;
  assign buffers_1_io_addrDebug = io_addrDebug_1; // @[DebugBufferWriters.scala 47:29]
  assign buffers_1_io_vmeOut_cmd_ready = io_vmeOut_1_cmd_ready; // @[DebugBufferWriters.scala 48:18]
  assign buffers_1_io_vmeOut_data_ready = io_vmeOut_1_data_ready; // @[DebugBufferWriters.scala 48:18]
  assign buffers_1_io_vmeOut_ack = io_vmeOut_1_ack; // @[DebugBufferWriters.scala 48:18]
  assign buffers_2_clock = clock;
  assign buffers_2_reset = reset;
  assign buffers_2_io_addrDebug = io_addrDebug_2; // @[DebugBufferWriters.scala 47:29]
  assign buffers_2_io_vmeOut_cmd_ready = io_vmeOut_2_cmd_ready; // @[DebugBufferWriters.scala 48:18]
  assign buffers_2_io_vmeOut_data_ready = io_vmeOut_2_data_ready; // @[DebugBufferWriters.scala 48:18]
  assign buffers_2_io_vmeOut_ack = io_vmeOut_2_ack; // @[DebugBufferWriters.scala 48:18]
endmodule
module DandelionDebugFPGAShell(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [15:0] io_host_aw_bits_addr,
  input  [12:0] io_host_aw_bits_id,
  input  [9:0]  io_host_aw_bits_user,
  input  [3:0]  io_host_aw_bits_len,
  input  [2:0]  io_host_aw_bits_size,
  input  [1:0]  io_host_aw_bits_burst,
  input  [1:0]  io_host_aw_bits_lock,
  input  [3:0]  io_host_aw_bits_cache,
  input  [2:0]  io_host_aw_bits_prot,
  input  [3:0]  io_host_aw_bits_qos,
  input  [3:0]  io_host_aw_bits_region,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [31:0] io_host_w_bits_data,
  input  [3:0]  io_host_w_bits_strb,
  input         io_host_w_bits_last,
  input  [12:0] io_host_w_bits_id,
  input  [9:0]  io_host_w_bits_user,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output [1:0]  io_host_b_bits_resp,
  output [12:0] io_host_b_bits_id,
  output [9:0]  io_host_b_bits_user,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [15:0] io_host_ar_bits_addr,
  input  [12:0] io_host_ar_bits_id,
  input  [9:0]  io_host_ar_bits_user,
  input  [3:0]  io_host_ar_bits_len,
  input  [2:0]  io_host_ar_bits_size,
  input  [1:0]  io_host_ar_bits_burst,
  input  [1:0]  io_host_ar_bits_lock,
  input  [3:0]  io_host_ar_bits_cache,
  input  [2:0]  io_host_ar_bits_prot,
  input  [3:0]  io_host_ar_bits_qos,
  input  [3:0]  io_host_ar_bits_region,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [31:0] io_host_r_bits_data,
  output [1:0]  io_host_r_bits_resp,
  output        io_host_r_bits_last,
  output [12:0] io_host_r_bits_id,
  output [9:0]  io_host_r_bits_user,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [15:0] io_mem_aw_bits_id,
  output [4:0]  io_mem_aw_bits_user,
  output [7:0]  io_mem_aw_bits_len,
  output [2:0]  io_mem_aw_bits_size,
  output [1:0]  io_mem_aw_bits_burst,
  output [1:0]  io_mem_aw_bits_lock,
  output [3:0]  io_mem_aw_bits_cache,
  output [2:0]  io_mem_aw_bits_prot,
  output [3:0]  io_mem_aw_bits_qos,
  output [3:0]  io_mem_aw_bits_region,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output [7:0]  io_mem_w_bits_strb,
  output        io_mem_w_bits_last,
  output [15:0] io_mem_w_bits_id,
  output [4:0]  io_mem_w_bits_user,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input  [1:0]  io_mem_b_bits_resp,
  input  [15:0] io_mem_b_bits_id,
  input  [4:0]  io_mem_b_bits_user,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [15:0] io_mem_ar_bits_id,
  output [4:0]  io_mem_ar_bits_user,
  output [7:0]  io_mem_ar_bits_len,
  output [2:0]  io_mem_ar_bits_size,
  output [1:0]  io_mem_ar_bits_burst,
  output [1:0]  io_mem_ar_bits_lock,
  output [3:0]  io_mem_ar_bits_cache,
  output [2:0]  io_mem_ar_bits_prot,
  output [3:0]  io_mem_ar_bits_qos,
  output [3:0]  io_mem_ar_bits_region,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input  [1:0]  io_mem_r_bits_resp,
  input         io_mem_r_bits_last,
  input  [15:0] io_mem_r_bits_id,
  input  [4:0]  io_mem_r_bits_user
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  dcr_clock; // @[DandelionShell.scala 817:19]
  wire  dcr_reset; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_aw_ready; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_aw_valid; // @[DandelionShell.scala 817:19]
  wire [15:0] dcr_io_host_aw_bits_addr; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_w_ready; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_w_valid; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_host_w_bits_data; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_b_ready; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_b_valid; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_ar_ready; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_ar_valid; // @[DandelionShell.scala 817:19]
  wire [15:0] dcr_io_host_ar_bits_addr; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_r_ready; // @[DandelionShell.scala 817:19]
  wire  dcr_io_host_r_valid; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_host_r_bits_data; // @[DandelionShell.scala 817:19]
  wire  dcr_io_dcr_launch; // @[DandelionShell.scala 817:19]
  wire  dcr_io_dcr_finish; // @[DandelionShell.scala 817:19]
  wire  dcr_io_dcr_ecnt_0_valid; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ecnt_0_bits; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ptrs_0; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ptrs_1; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ptrs_2; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ptrs_3; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ptrs_4; // @[DandelionShell.scala 817:19]
  wire [31:0] dcr_io_dcr_ptrs_5; // @[DandelionShell.scala 817:19]
  wire  dmem_clock; // @[DandelionShell.scala 818:20]
  wire  dmem_reset; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_aw_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_aw_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_mem_aw_bits_addr; // @[DandelionShell.scala 818:20]
  wire [7:0] dmem_io_mem_aw_bits_len; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_w_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_w_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_mem_w_bits_data; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_w_bits_last; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_b_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_b_valid; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_ar_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_ar_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_mem_ar_bits_addr; // @[DandelionShell.scala 818:20]
  wire [7:0] dmem_io_mem_ar_bits_len; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_r_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_r_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_mem_r_bits_data; // @[DandelionShell.scala 818:20]
  wire  dmem_io_mem_r_bits_last; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_rd_0_cmd_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_rd_0_cmd_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_dme_rd_0_cmd_bits_addr; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_rd_0_data_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_rd_0_data_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_dme_rd_0_data_bits; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_0_cmd_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_0_cmd_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_dme_wr_0_cmd_bits_addr; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_0_data_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_0_data_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_dme_wr_0_data_bits; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_0_ack; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_1_cmd_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_1_cmd_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_dme_wr_1_cmd_bits_addr; // @[DandelionShell.scala 818:20]
  wire [7:0] dmem_io_dme_wr_1_cmd_bits_len; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_1_data_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_1_data_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_dme_wr_1_data_bits; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_1_ack; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_2_cmd_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_2_cmd_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_dme_wr_2_cmd_bits_addr; // @[DandelionShell.scala 818:20]
  wire [7:0] dmem_io_dme_wr_2_cmd_bits_len; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_2_data_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_2_data_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_dme_wr_2_data_bits; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_2_ack; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_3_cmd_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_3_cmd_valid; // @[DandelionShell.scala 818:20]
  wire [31:0] dmem_io_dme_wr_3_cmd_bits_addr; // @[DandelionShell.scala 818:20]
  wire [7:0] dmem_io_dme_wr_3_cmd_bits_len; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_3_data_ready; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_3_data_valid; // @[DandelionShell.scala 818:20]
  wire [63:0] dmem_io_dme_wr_3_data_bits; // @[DandelionShell.scala 818:20]
  wire  dmem_io_dme_wr_3_ack; // @[DandelionShell.scala 818:20]
  wire  cache_clock; // @[DandelionShell.scala 819:21]
  wire  cache_reset; // @[DandelionShell.scala 819:21]
  wire  cache_io_cpu_flush; // @[DandelionShell.scala 819:21]
  wire  cache_io_cpu_flush_done; // @[DandelionShell.scala 819:21]
  wire  cache_io_cpu_req_ready; // @[DandelionShell.scala 819:21]
  wire  cache_io_cpu_req_valid; // @[DandelionShell.scala 819:21]
  wire [63:0] cache_io_cpu_req_bits_addr; // @[DandelionShell.scala 819:21]
  wire [63:0] cache_io_cpu_req_bits_data; // @[DandelionShell.scala 819:21]
  wire [7:0] cache_io_cpu_req_bits_mask; // @[DandelionShell.scala 819:21]
  wire [7:0] cache_io_cpu_req_bits_tag; // @[DandelionShell.scala 819:21]
  wire  cache_io_cpu_resp_valid; // @[DandelionShell.scala 819:21]
  wire [63:0] cache_io_cpu_resp_bits_data; // @[DandelionShell.scala 819:21]
  wire [7:0] cache_io_cpu_resp_bits_tag; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_rd_cmd_ready; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_rd_cmd_valid; // @[DandelionShell.scala 819:21]
  wire [31:0] cache_io_mem_rd_cmd_bits_addr; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_rd_data_ready; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_rd_data_valid; // @[DandelionShell.scala 819:21]
  wire [63:0] cache_io_mem_rd_data_bits; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_wr_cmd_ready; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_wr_cmd_valid; // @[DandelionShell.scala 819:21]
  wire [31:0] cache_io_mem_wr_cmd_bits_addr; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_wr_data_ready; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_wr_data_valid; // @[DandelionShell.scala 819:21]
  wire [63:0] cache_io_mem_wr_data_bits; // @[DandelionShell.scala 819:21]
  wire  cache_io_mem_wr_ack; // @[DandelionShell.scala 819:21]
  wire  accel_clock; // @[DandelionShell.scala 822:21]
  wire  accel_reset; // @[DandelionShell.scala 822:21]
  wire  accel_io_in_ready; // @[DandelionShell.scala 822:21]
  wire  accel_io_in_valid; // @[DandelionShell.scala 822:21]
  wire [31:0] accel_io_in_bits_dataPtrs_field2_data; // @[DandelionShell.scala 822:21]
  wire [31:0] accel_io_in_bits_dataPtrs_field1_data; // @[DandelionShell.scala 822:21]
  wire [31:0] accel_io_in_bits_dataPtrs_field0_data; // @[DandelionShell.scala 822:21]
  wire  accel_io_MemResp_valid; // @[DandelionShell.scala 822:21]
  wire [63:0] accel_io_MemResp_bits_data; // @[DandelionShell.scala 822:21]
  wire [7:0] accel_io_MemResp_bits_tag; // @[DandelionShell.scala 822:21]
  wire  accel_io_MemReq_ready; // @[DandelionShell.scala 822:21]
  wire  accel_io_MemReq_valid; // @[DandelionShell.scala 822:21]
  wire [63:0] accel_io_MemReq_bits_addr; // @[DandelionShell.scala 822:21]
  wire [63:0] accel_io_MemReq_bits_data; // @[DandelionShell.scala 822:21]
  wire [7:0] accel_io_MemReq_bits_mask; // @[DandelionShell.scala 822:21]
  wire [7:0] accel_io_MemReq_bits_tag; // @[DandelionShell.scala 822:21]
  wire  accel_io_out_ready; // @[DandelionShell.scala 822:21]
  wire  accel_io_out_valid; // @[DandelionShell.scala 822:21]
  wire  debug_module_clock; // @[DandelionShell.scala 824:50]
  wire  debug_module_reset; // @[DandelionShell.scala 824:50]
  wire [31:0] debug_module_io_addrDebug_0; // @[DandelionShell.scala 824:50]
  wire [31:0] debug_module_io_addrDebug_1; // @[DandelionShell.scala 824:50]
  wire [31:0] debug_module_io_addrDebug_2; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_0_cmd_ready; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_0_cmd_valid; // @[DandelionShell.scala 824:50]
  wire [31:0] debug_module_io_vmeOut_0_cmd_bits_addr; // @[DandelionShell.scala 824:50]
  wire [7:0] debug_module_io_vmeOut_0_cmd_bits_len; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_0_data_ready; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_0_data_valid; // @[DandelionShell.scala 824:50]
  wire [63:0] debug_module_io_vmeOut_0_data_bits; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_0_ack; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_1_cmd_ready; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_1_cmd_valid; // @[DandelionShell.scala 824:50]
  wire [31:0] debug_module_io_vmeOut_1_cmd_bits_addr; // @[DandelionShell.scala 824:50]
  wire [7:0] debug_module_io_vmeOut_1_cmd_bits_len; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_1_data_ready; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_1_data_valid; // @[DandelionShell.scala 824:50]
  wire [63:0] debug_module_io_vmeOut_1_data_bits; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_1_ack; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_2_cmd_ready; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_2_cmd_valid; // @[DandelionShell.scala 824:50]
  wire [31:0] debug_module_io_vmeOut_2_cmd_bits_addr; // @[DandelionShell.scala 824:50]
  wire [7:0] debug_module_io_vmeOut_2_cmd_bits_len; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_2_data_ready; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_2_data_valid; // @[DandelionShell.scala 824:50]
  wire [63:0] debug_module_io_vmeOut_2_data_bits; // @[DandelionShell.scala 824:50]
  wire  debug_module_io_vmeOut_2_ack; // @[DandelionShell.scala 824:50]
  reg [1:0] state; // @[DandelionShell.scala 843:22]
  reg [31:0] cycles; // @[DandelionShell.scala 844:23]
  wire  _T = state == 2'h0; // @[DandelionShell.scala 849:14]
  wire  _T_1 = state != 2'h2; // @[DandelionShell.scala 851:20]
  wire [31:0] _T_3 = cycles + 32'h1; // @[DandelionShell.scala 852:22]
  reg [63:0] ptrs_0; // @[Reg.scala 27:20]
  reg [63:0] ptrs_1; // @[Reg.scala 27:20]
  reg [63:0] ptrs_2; // @[Reg.scala 27:20]
  reg [63:0] ptrs_3; // @[Reg.scala 27:20]
  reg [63:0] ptrs_4; // @[Reg.scala 27:20]
  reg [63:0] ptrs_5; // @[Reg.scala 27:20]
  wire  _T_14 = state == 2'h2; // @[DandelionShell.scala 900:31]
  reg  dme_ack_0; // @[DandelionShell.scala 911:46]
  reg  dme_ack_1; // @[DandelionShell.scala 911:46]
  reg  dme_ack_2; // @[DandelionShell.scala 911:46]
  wire  _GEN_8 = dmem_io_dme_wr_1_ack | dme_ack_0; // @[DandelionShell.scala 913:37]
  wire  _GEN_9 = dmem_io_dme_wr_2_ack | dme_ack_1; // @[DandelionShell.scala 913:37]
  wire  _GEN_10 = dmem_io_dme_wr_3_ack | dme_ack_2; // @[DandelionShell.scala 913:37]
  reg  cache_done; // @[DandelionShell.scala 926:27]
  wire  _GEN_11 = cache_io_cpu_flush_done | cache_done; // @[DandelionShell.scala 928:35]
  wire  _T_17 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = ~reset; // @[DandelionShell.scala 936:15]
  wire  _T_38 = accel_io_in_ready & accel_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_14 = dcr_io_dcr_launch; // @[DandelionShell.scala 935:31]
  wire  _T_39 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_40 = accel_io_out_ready & accel_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_41 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_42 = dme_ack_0 & dme_ack_1; // @[DandelionShell.scala 922:32]
  wire  _T_43 = _T_42 & dme_ack_2; // @[DandelionShell.scala 922:32]
  wire  _T_44 = cache_done & _T_43; // @[DandelionShell.scala 957:23]
  wire  _T_45 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire  _GEN_23 = _T_17 & dcr_io_dcr_launch; // @[DandelionShell.scala 936:15]
  DCR dcr ( // @[DandelionShell.scala 817:19]
    .clock(dcr_clock),
    .reset(dcr_reset),
    .io_host_aw_ready(dcr_io_host_aw_ready),
    .io_host_aw_valid(dcr_io_host_aw_valid),
    .io_host_aw_bits_addr(dcr_io_host_aw_bits_addr),
    .io_host_w_ready(dcr_io_host_w_ready),
    .io_host_w_valid(dcr_io_host_w_valid),
    .io_host_w_bits_data(dcr_io_host_w_bits_data),
    .io_host_b_ready(dcr_io_host_b_ready),
    .io_host_b_valid(dcr_io_host_b_valid),
    .io_host_ar_ready(dcr_io_host_ar_ready),
    .io_host_ar_valid(dcr_io_host_ar_valid),
    .io_host_ar_bits_addr(dcr_io_host_ar_bits_addr),
    .io_host_r_ready(dcr_io_host_r_ready),
    .io_host_r_valid(dcr_io_host_r_valid),
    .io_host_r_bits_data(dcr_io_host_r_bits_data),
    .io_dcr_launch(dcr_io_dcr_launch),
    .io_dcr_finish(dcr_io_dcr_finish),
    .io_dcr_ecnt_0_valid(dcr_io_dcr_ecnt_0_valid),
    .io_dcr_ecnt_0_bits(dcr_io_dcr_ecnt_0_bits),
    .io_dcr_ptrs_0(dcr_io_dcr_ptrs_0),
    .io_dcr_ptrs_1(dcr_io_dcr_ptrs_1),
    .io_dcr_ptrs_2(dcr_io_dcr_ptrs_2),
    .io_dcr_ptrs_3(dcr_io_dcr_ptrs_3),
    .io_dcr_ptrs_4(dcr_io_dcr_ptrs_4),
    .io_dcr_ptrs_5(dcr_io_dcr_ptrs_5)
  );
  DME dmem ( // @[DandelionShell.scala 818:20]
    .clock(dmem_clock),
    .reset(dmem_reset),
    .io_mem_aw_ready(dmem_io_mem_aw_ready),
    .io_mem_aw_valid(dmem_io_mem_aw_valid),
    .io_mem_aw_bits_addr(dmem_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(dmem_io_mem_aw_bits_len),
    .io_mem_w_ready(dmem_io_mem_w_ready),
    .io_mem_w_valid(dmem_io_mem_w_valid),
    .io_mem_w_bits_data(dmem_io_mem_w_bits_data),
    .io_mem_w_bits_last(dmem_io_mem_w_bits_last),
    .io_mem_b_ready(dmem_io_mem_b_ready),
    .io_mem_b_valid(dmem_io_mem_b_valid),
    .io_mem_ar_ready(dmem_io_mem_ar_ready),
    .io_mem_ar_valid(dmem_io_mem_ar_valid),
    .io_mem_ar_bits_addr(dmem_io_mem_ar_bits_addr),
    .io_mem_ar_bits_len(dmem_io_mem_ar_bits_len),
    .io_mem_r_ready(dmem_io_mem_r_ready),
    .io_mem_r_valid(dmem_io_mem_r_valid),
    .io_mem_r_bits_data(dmem_io_mem_r_bits_data),
    .io_mem_r_bits_last(dmem_io_mem_r_bits_last),
    .io_dme_rd_0_cmd_ready(dmem_io_dme_rd_0_cmd_ready),
    .io_dme_rd_0_cmd_valid(dmem_io_dme_rd_0_cmd_valid),
    .io_dme_rd_0_cmd_bits_addr(dmem_io_dme_rd_0_cmd_bits_addr),
    .io_dme_rd_0_data_ready(dmem_io_dme_rd_0_data_ready),
    .io_dme_rd_0_data_valid(dmem_io_dme_rd_0_data_valid),
    .io_dme_rd_0_data_bits(dmem_io_dme_rd_0_data_bits),
    .io_dme_wr_0_cmd_ready(dmem_io_dme_wr_0_cmd_ready),
    .io_dme_wr_0_cmd_valid(dmem_io_dme_wr_0_cmd_valid),
    .io_dme_wr_0_cmd_bits_addr(dmem_io_dme_wr_0_cmd_bits_addr),
    .io_dme_wr_0_data_ready(dmem_io_dme_wr_0_data_ready),
    .io_dme_wr_0_data_valid(dmem_io_dme_wr_0_data_valid),
    .io_dme_wr_0_data_bits(dmem_io_dme_wr_0_data_bits),
    .io_dme_wr_0_ack(dmem_io_dme_wr_0_ack),
    .io_dme_wr_1_cmd_ready(dmem_io_dme_wr_1_cmd_ready),
    .io_dme_wr_1_cmd_valid(dmem_io_dme_wr_1_cmd_valid),
    .io_dme_wr_1_cmd_bits_addr(dmem_io_dme_wr_1_cmd_bits_addr),
    .io_dme_wr_1_cmd_bits_len(dmem_io_dme_wr_1_cmd_bits_len),
    .io_dme_wr_1_data_ready(dmem_io_dme_wr_1_data_ready),
    .io_dme_wr_1_data_valid(dmem_io_dme_wr_1_data_valid),
    .io_dme_wr_1_data_bits(dmem_io_dme_wr_1_data_bits),
    .io_dme_wr_1_ack(dmem_io_dme_wr_1_ack),
    .io_dme_wr_2_cmd_ready(dmem_io_dme_wr_2_cmd_ready),
    .io_dme_wr_2_cmd_valid(dmem_io_dme_wr_2_cmd_valid),
    .io_dme_wr_2_cmd_bits_addr(dmem_io_dme_wr_2_cmd_bits_addr),
    .io_dme_wr_2_cmd_bits_len(dmem_io_dme_wr_2_cmd_bits_len),
    .io_dme_wr_2_data_ready(dmem_io_dme_wr_2_data_ready),
    .io_dme_wr_2_data_valid(dmem_io_dme_wr_2_data_valid),
    .io_dme_wr_2_data_bits(dmem_io_dme_wr_2_data_bits),
    .io_dme_wr_2_ack(dmem_io_dme_wr_2_ack),
    .io_dme_wr_3_cmd_ready(dmem_io_dme_wr_3_cmd_ready),
    .io_dme_wr_3_cmd_valid(dmem_io_dme_wr_3_cmd_valid),
    .io_dme_wr_3_cmd_bits_addr(dmem_io_dme_wr_3_cmd_bits_addr),
    .io_dme_wr_3_cmd_bits_len(dmem_io_dme_wr_3_cmd_bits_len),
    .io_dme_wr_3_data_ready(dmem_io_dme_wr_3_data_ready),
    .io_dme_wr_3_data_valid(dmem_io_dme_wr_3_data_valid),
    .io_dme_wr_3_data_bits(dmem_io_dme_wr_3_data_bits),
    .io_dme_wr_3_ack(dmem_io_dme_wr_3_ack)
  );
  DMECache cache ( // @[DandelionShell.scala 819:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .io_cpu_flush(cache_io_cpu_flush),
    .io_cpu_flush_done(cache_io_cpu_flush_done),
    .io_cpu_req_ready(cache_io_cpu_req_ready),
    .io_cpu_req_valid(cache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(cache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(cache_io_cpu_req_bits_data),
    .io_cpu_req_bits_mask(cache_io_cpu_req_bits_mask),
    .io_cpu_req_bits_tag(cache_io_cpu_req_bits_tag),
    .io_cpu_resp_valid(cache_io_cpu_resp_valid),
    .io_cpu_resp_bits_data(cache_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_tag(cache_io_cpu_resp_bits_tag),
    .io_mem_rd_cmd_ready(cache_io_mem_rd_cmd_ready),
    .io_mem_rd_cmd_valid(cache_io_mem_rd_cmd_valid),
    .io_mem_rd_cmd_bits_addr(cache_io_mem_rd_cmd_bits_addr),
    .io_mem_rd_data_ready(cache_io_mem_rd_data_ready),
    .io_mem_rd_data_valid(cache_io_mem_rd_data_valid),
    .io_mem_rd_data_bits(cache_io_mem_rd_data_bits),
    .io_mem_wr_cmd_ready(cache_io_mem_wr_cmd_ready),
    .io_mem_wr_cmd_valid(cache_io_mem_wr_cmd_valid),
    .io_mem_wr_cmd_bits_addr(cache_io_mem_wr_cmd_bits_addr),
    .io_mem_wr_data_ready(cache_io_mem_wr_data_ready),
    .io_mem_wr_data_valid(cache_io_mem_wr_data_valid),
    .io_mem_wr_data_bits(cache_io_mem_wr_data_bits),
    .io_mem_wr_ack(cache_io_mem_wr_ack)
  );
  bbgemmDF accel ( // @[DandelionShell.scala 822:21]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_in_ready(accel_io_in_ready),
    .io_in_valid(accel_io_in_valid),
    .io_in_bits_dataPtrs_field2_data(accel_io_in_bits_dataPtrs_field2_data),
    .io_in_bits_dataPtrs_field1_data(accel_io_in_bits_dataPtrs_field1_data),
    .io_in_bits_dataPtrs_field0_data(accel_io_in_bits_dataPtrs_field0_data),
    .io_MemResp_valid(accel_io_MemResp_valid),
    .io_MemResp_bits_data(accel_io_MemResp_bits_data),
    .io_MemResp_bits_tag(accel_io_MemResp_bits_tag),
    .io_MemReq_ready(accel_io_MemReq_ready),
    .io_MemReq_valid(accel_io_MemReq_valid),
    .io_MemReq_bits_addr(accel_io_MemReq_bits_addr),
    .io_MemReq_bits_data(accel_io_MemReq_bits_data),
    .io_MemReq_bits_mask(accel_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(accel_io_MemReq_bits_tag),
    .io_out_ready(accel_io_out_ready),
    .io_out_valid(accel_io_out_valid)
  );
  DebugBufferWriters debug_module ( // @[DandelionShell.scala 824:50]
    .clock(debug_module_clock),
    .reset(debug_module_reset),
    .io_addrDebug_0(debug_module_io_addrDebug_0),
    .io_addrDebug_1(debug_module_io_addrDebug_1),
    .io_addrDebug_2(debug_module_io_addrDebug_2),
    .io_vmeOut_0_cmd_ready(debug_module_io_vmeOut_0_cmd_ready),
    .io_vmeOut_0_cmd_valid(debug_module_io_vmeOut_0_cmd_valid),
    .io_vmeOut_0_cmd_bits_addr(debug_module_io_vmeOut_0_cmd_bits_addr),
    .io_vmeOut_0_cmd_bits_len(debug_module_io_vmeOut_0_cmd_bits_len),
    .io_vmeOut_0_data_ready(debug_module_io_vmeOut_0_data_ready),
    .io_vmeOut_0_data_valid(debug_module_io_vmeOut_0_data_valid),
    .io_vmeOut_0_data_bits(debug_module_io_vmeOut_0_data_bits),
    .io_vmeOut_0_ack(debug_module_io_vmeOut_0_ack),
    .io_vmeOut_1_cmd_ready(debug_module_io_vmeOut_1_cmd_ready),
    .io_vmeOut_1_cmd_valid(debug_module_io_vmeOut_1_cmd_valid),
    .io_vmeOut_1_cmd_bits_addr(debug_module_io_vmeOut_1_cmd_bits_addr),
    .io_vmeOut_1_cmd_bits_len(debug_module_io_vmeOut_1_cmd_bits_len),
    .io_vmeOut_1_data_ready(debug_module_io_vmeOut_1_data_ready),
    .io_vmeOut_1_data_valid(debug_module_io_vmeOut_1_data_valid),
    .io_vmeOut_1_data_bits(debug_module_io_vmeOut_1_data_bits),
    .io_vmeOut_1_ack(debug_module_io_vmeOut_1_ack),
    .io_vmeOut_2_cmd_ready(debug_module_io_vmeOut_2_cmd_ready),
    .io_vmeOut_2_cmd_valid(debug_module_io_vmeOut_2_cmd_valid),
    .io_vmeOut_2_cmd_bits_addr(debug_module_io_vmeOut_2_cmd_bits_addr),
    .io_vmeOut_2_cmd_bits_len(debug_module_io_vmeOut_2_cmd_bits_len),
    .io_vmeOut_2_data_ready(debug_module_io_vmeOut_2_data_ready),
    .io_vmeOut_2_data_valid(debug_module_io_vmeOut_2_data_valid),
    .io_vmeOut_2_data_bits(debug_module_io_vmeOut_2_data_bits),
    .io_vmeOut_2_ack(debug_module_io_vmeOut_2_ack)
  );
  assign io_host_aw_ready = dcr_io_host_aw_ready; // @[DandelionShell.scala 970:11]
  assign io_host_w_ready = dcr_io_host_w_ready; // @[DandelionShell.scala 970:11]
  assign io_host_b_valid = dcr_io_host_b_valid; // @[DandelionShell.scala 970:11]
  assign io_host_b_bits_resp = 2'h0; // @[DandelionShell.scala 970:11]
  assign io_host_b_bits_id = io_host_w_bits_id; // @[DandelionShell.scala 973:21]
  assign io_host_b_bits_user = 10'h0;
  assign io_host_ar_ready = dcr_io_host_ar_ready; // @[DandelionShell.scala 970:11]
  assign io_host_r_valid = dcr_io_host_r_valid; // @[DandelionShell.scala 970:11]
  assign io_host_r_bits_data = dcr_io_host_r_bits_data; // @[DandelionShell.scala 970:11]
  assign io_host_r_bits_resp = 2'h0; // @[DandelionShell.scala 970:11]
  assign io_host_r_bits_last = 1'h1; // @[DandelionShell.scala 978:23]
  assign io_host_r_bits_id = io_host_ar_bits_id; // @[DandelionShell.scala 974:21]
  assign io_host_r_bits_user = 10'h0;
  assign io_mem_aw_valid = dmem_io_mem_aw_valid; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_addr = dmem_io_mem_aw_bits_addr; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_id = 16'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_user = 5'h1; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_len = dmem_io_mem_aw_bits_len; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_size = 3'h3; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_burst = 2'h1; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_lock = 2'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_cache = 4'hf; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_prot = 3'h4; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_qos = 4'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_aw_bits_region = 4'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_w_valid = dmem_io_mem_w_valid; // @[DandelionShell.scala 969:10]
  assign io_mem_w_bits_data = dmem_io_mem_w_bits_data; // @[DandelionShell.scala 969:10]
  assign io_mem_w_bits_strb = 8'hff; // @[DandelionShell.scala 969:10]
  assign io_mem_w_bits_last = dmem_io_mem_w_bits_last; // @[DandelionShell.scala 969:10]
  assign io_mem_w_bits_id = 16'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_w_bits_user = 5'h1; // @[DandelionShell.scala 969:10]
  assign io_mem_b_ready = dmem_io_mem_b_ready; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_valid = dmem_io_mem_ar_valid; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_addr = dmem_io_mem_ar_bits_addr; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_id = 16'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_user = 5'h1; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_len = dmem_io_mem_ar_bits_len; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_size = 3'h3; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_burst = 2'h1; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_lock = 2'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_cache = 4'hf; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_prot = 3'h4; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_qos = 4'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_ar_bits_region = 4'h0; // @[DandelionShell.scala 969:10]
  assign io_mem_r_ready = dmem_io_mem_r_ready; // @[DandelionShell.scala 969:10]
  assign dcr_clock = clock;
  assign dcr_reset = reset;
  assign dcr_io_host_aw_valid = io_host_aw_valid; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_aw_bits_addr = io_host_aw_bits_addr; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_w_valid = io_host_w_valid; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_w_bits_data = io_host_w_bits_data; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_b_ready = io_host_b_ready; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_ar_valid = io_host_ar_valid; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_ar_bits_addr = io_host_ar_bits_addr; // @[DandelionShell.scala 970:11]
  assign dcr_io_host_r_ready = io_host_r_ready; // @[DandelionShell.scala 970:11]
  assign dcr_io_dcr_finish = state == 2'h3; // @[DandelionShell.scala 967:21]
  assign dcr_io_dcr_ecnt_0_valid = state == 2'h3; // @[DandelionShell.scala 859:28]
  assign dcr_io_dcr_ecnt_0_bits = cycles; // @[DandelionShell.scala 860:27]
  assign dmem_clock = clock;
  assign dmem_reset = reset;
  assign dmem_io_mem_aw_ready = io_mem_aw_ready; // @[DandelionShell.scala 969:10]
  assign dmem_io_mem_w_ready = io_mem_w_ready; // @[DandelionShell.scala 969:10]
  assign dmem_io_mem_b_valid = io_mem_b_valid; // @[DandelionShell.scala 969:10]
  assign dmem_io_mem_ar_ready = io_mem_ar_ready; // @[DandelionShell.scala 969:10]
  assign dmem_io_mem_r_valid = io_mem_r_valid; // @[DandelionShell.scala 969:10]
  assign dmem_io_mem_r_bits_data = io_mem_r_bits_data; // @[DandelionShell.scala 969:10]
  assign dmem_io_mem_r_bits_last = io_mem_r_bits_last; // @[DandelionShell.scala 969:10]
  assign dmem_io_dme_rd_0_cmd_valid = cache_io_mem_rd_cmd_valid; // @[DandelionShell.scala 833:21]
  assign dmem_io_dme_rd_0_cmd_bits_addr = cache_io_mem_rd_cmd_bits_addr; // @[DandelionShell.scala 833:21]
  assign dmem_io_dme_rd_0_data_ready = cache_io_mem_rd_data_ready; // @[DandelionShell.scala 833:21]
  assign dmem_io_dme_wr_0_cmd_valid = cache_io_mem_wr_cmd_valid; // @[DandelionShell.scala 834:21]
  assign dmem_io_dme_wr_0_cmd_bits_addr = cache_io_mem_wr_cmd_bits_addr; // @[DandelionShell.scala 834:21]
  assign dmem_io_dme_wr_0_data_valid = cache_io_mem_wr_data_valid; // @[DandelionShell.scala 834:21]
  assign dmem_io_dme_wr_0_data_bits = cache_io_mem_wr_data_bits; // @[DandelionShell.scala 834:21]
  assign dmem_io_dme_wr_1_cmd_valid = debug_module_io_vmeOut_0_cmd_valid; // @[DandelionShell.scala 904:37]
  assign dmem_io_dme_wr_1_cmd_bits_addr = debug_module_io_vmeOut_0_cmd_bits_addr; // @[DandelionShell.scala 903:36]
  assign dmem_io_dme_wr_1_cmd_bits_len = debug_module_io_vmeOut_0_cmd_bits_len; // @[DandelionShell.scala 903:36]
  assign dmem_io_dme_wr_1_data_valid = debug_module_io_vmeOut_0_data_valid; // @[DandelionShell.scala 907:32]
  assign dmem_io_dme_wr_1_data_bits = debug_module_io_vmeOut_0_data_bits; // @[DandelionShell.scala 907:32]
  assign dmem_io_dme_wr_2_cmd_valid = debug_module_io_vmeOut_1_cmd_valid; // @[DandelionShell.scala 904:37]
  assign dmem_io_dme_wr_2_cmd_bits_addr = debug_module_io_vmeOut_1_cmd_bits_addr; // @[DandelionShell.scala 903:36]
  assign dmem_io_dme_wr_2_cmd_bits_len = debug_module_io_vmeOut_1_cmd_bits_len; // @[DandelionShell.scala 903:36]
  assign dmem_io_dme_wr_2_data_valid = debug_module_io_vmeOut_1_data_valid; // @[DandelionShell.scala 907:32]
  assign dmem_io_dme_wr_2_data_bits = debug_module_io_vmeOut_1_data_bits; // @[DandelionShell.scala 907:32]
  assign dmem_io_dme_wr_3_cmd_valid = debug_module_io_vmeOut_2_cmd_valid; // @[DandelionShell.scala 904:37]
  assign dmem_io_dme_wr_3_cmd_bits_addr = debug_module_io_vmeOut_2_cmd_bits_addr; // @[DandelionShell.scala 903:36]
  assign dmem_io_dme_wr_3_cmd_bits_len = debug_module_io_vmeOut_2_cmd_bits_len; // @[DandelionShell.scala 903:36]
  assign dmem_io_dme_wr_3_data_valid = debug_module_io_vmeOut_2_data_valid; // @[DandelionShell.scala 907:32]
  assign dmem_io_dme_wr_3_data_bits = debug_module_io_vmeOut_2_data_bits; // @[DandelionShell.scala 907:32]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_io_cpu_flush = state == 2'h2; // @[DandelionShell.scala 900:22]
  assign cache_io_cpu_req_valid = accel_io_MemReq_valid; // @[DandelionShell.scala 826:20]
  assign cache_io_cpu_req_bits_addr = accel_io_MemReq_bits_addr; // @[DandelionShell.scala 826:20]
  assign cache_io_cpu_req_bits_data = accel_io_MemReq_bits_data; // @[DandelionShell.scala 826:20]
  assign cache_io_cpu_req_bits_mask = accel_io_MemReq_bits_mask; // @[DandelionShell.scala 826:20]
  assign cache_io_cpu_req_bits_tag = accel_io_MemReq_bits_tag; // @[DandelionShell.scala 826:20]
  assign cache_io_mem_rd_cmd_ready = dmem_io_dme_rd_0_cmd_ready; // @[DandelionShell.scala 833:21]
  assign cache_io_mem_rd_data_valid = dmem_io_dme_rd_0_data_valid; // @[DandelionShell.scala 833:21]
  assign cache_io_mem_rd_data_bits = dmem_io_dme_rd_0_data_bits; // @[DandelionShell.scala 833:21]
  assign cache_io_mem_wr_cmd_ready = dmem_io_dme_wr_0_cmd_ready; // @[DandelionShell.scala 834:21]
  assign cache_io_mem_wr_data_ready = dmem_io_dme_wr_0_data_ready; // @[DandelionShell.scala 834:21]
  assign cache_io_mem_wr_ack = dmem_io_dme_wr_0_ack; // @[DandelionShell.scala 834:21]
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign accel_io_in_valid = _T_17 & _GEN_14; // @[DandelionShell.scala 897:21 DandelionShell.scala 945:27]
  assign accel_io_in_bits_dataPtrs_field2_data = ptrs_2[31:0]; // @[DandelionShell.scala 879:45]
  assign accel_io_in_bits_dataPtrs_field1_data = ptrs_1[31:0]; // @[DandelionShell.scala 879:45]
  assign accel_io_in_bits_dataPtrs_field0_data = ptrs_0[31:0]; // @[DandelionShell.scala 879:45]
  assign accel_io_MemResp_valid = cache_io_cpu_resp_valid; // @[DandelionShell.scala 827:20]
  assign accel_io_MemResp_bits_data = cache_io_cpu_resp_bits_data; // @[DandelionShell.scala 827:20]
  assign accel_io_MemResp_bits_tag = cache_io_cpu_resp_bits_tag; // @[DandelionShell.scala 827:20]
  assign accel_io_MemReq_ready = cache_io_cpu_req_ready; // @[DandelionShell.scala 826:20]
  assign accel_io_out_ready = state == 2'h1; // @[DandelionShell.scala 898:22]
  assign debug_module_clock = clock;
  assign debug_module_reset = reset;
  assign debug_module_io_addrDebug_0 = dcr_io_dcr_ptrs_3; // @[DandelionShell.scala 886:38]
  assign debug_module_io_addrDebug_1 = dcr_io_dcr_ptrs_4; // @[DandelionShell.scala 886:38]
  assign debug_module_io_addrDebug_2 = dcr_io_dcr_ptrs_5; // @[DandelionShell.scala 886:38]
  assign debug_module_io_vmeOut_0_cmd_ready = dmem_io_dme_wr_1_cmd_ready; // @[DandelionShell.scala 905:45]
  assign debug_module_io_vmeOut_0_data_ready = dmem_io_dme_wr_1_data_ready; // @[DandelionShell.scala 907:32]
  assign debug_module_io_vmeOut_0_ack = dmem_io_dme_wr_1_ack; // @[DandelionShell.scala 908:39]
  assign debug_module_io_vmeOut_1_cmd_ready = dmem_io_dme_wr_2_cmd_ready; // @[DandelionShell.scala 905:45]
  assign debug_module_io_vmeOut_1_data_ready = dmem_io_dme_wr_2_data_ready; // @[DandelionShell.scala 907:32]
  assign debug_module_io_vmeOut_1_ack = dmem_io_dme_wr_2_ack; // @[DandelionShell.scala 908:39]
  assign debug_module_io_vmeOut_2_cmd_ready = dmem_io_dme_wr_3_cmd_ready; // @[DandelionShell.scala 905:45]
  assign debug_module_io_vmeOut_2_data_ready = dmem_io_dme_wr_3_data_ready; // @[DandelionShell.scala 907:32]
  assign debug_module_io_vmeOut_2_ack = dmem_io_dme_wr_3_ack; // @[DandelionShell.scala 908:39]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  cycles = _RAND_1[31:0];
  _RAND_2 = {2{`RANDOM}};
  ptrs_0 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  ptrs_1 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  ptrs_2 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ptrs_3 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  ptrs_4 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  ptrs_5 = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  dme_ack_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dme_ack_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  dme_ack_2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cache_done = _RAND_11[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_17) begin
      if (dcr_io_dcr_launch) begin
        if (_T_38) begin
          state <= 2'h1;
        end
      end
    end else if (_T_39) begin
      if (_T_40) begin
        state <= 2'h2;
      end
    end else if (_T_41) begin
      if (_T_44) begin
        state <= 2'h3;
      end
    end else if (_T_45) begin
      state <= 2'h0;
    end
    if (reset) begin
      cycles <= 32'h0;
    end else if (_T) begin
      cycles <= 32'h0;
    end else if (_T_1) begin
      cycles <= _T_3;
    end
    if (reset) begin
      ptrs_0 <= 64'h0;
    end else if (_T) begin
      ptrs_0 <= {{32'd0}, dcr_io_dcr_ptrs_0};
    end
    if (reset) begin
      ptrs_1 <= 64'h0;
    end else if (_T) begin
      ptrs_1 <= {{32'd0}, dcr_io_dcr_ptrs_1};
    end
    if (reset) begin
      ptrs_2 <= 64'h0;
    end else if (_T) begin
      ptrs_2 <= {{32'd0}, dcr_io_dcr_ptrs_2};
    end
    if (reset) begin
      ptrs_3 <= 64'h0;
    end else if (_T) begin
      ptrs_3 <= {{32'd0}, dcr_io_dcr_ptrs_3};
    end
    if (reset) begin
      ptrs_4 <= 64'h0;
    end else if (_T) begin
      ptrs_4 <= {{32'd0}, dcr_io_dcr_ptrs_4};
    end
    if (reset) begin
      ptrs_5 <= 64'h0;
    end else if (_T) begin
      ptrs_5 <= {{32'd0}, dcr_io_dcr_ptrs_5};
    end
    if (reset) begin
      dme_ack_0 <= 1'h0;
    end else begin
      dme_ack_0 <= _GEN_8;
    end
    if (reset) begin
      dme_ack_1 <= 1'h0;
    end else begin
      dme_ack_1 <= _GEN_9;
    end
    if (reset) begin
      dme_ack_2 <= 1'h0;
    end else begin
      dme_ack_2 <= _GEN_10;
    end
    if (reset) begin
      cache_done <= 1'h0;
    end else if (_T_14) begin
      cache_done <= _GEN_11;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"Ptrs: "); // @[DandelionShell.scala 936:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"ptr(0): 0x%x, ",ptrs_0); // @[DandelionShell.scala 937:46]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"ptr(1): 0x%x, ",ptrs_1); // @[DandelionShell.scala 937:46]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"ptr(2): 0x%x, ",ptrs_2); // @[DandelionShell.scala 937:46]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"ptr(3): 0x%x, ",ptrs_3); // @[DandelionShell.scala 937:46]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"ptr(4): 0x%x, ",ptrs_4); // @[DandelionShell.scala 937:46]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"ptr(5): 0x%x, ",ptrs_5); // @[DandelionShell.scala 937:46]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"\nVals: "); // @[DandelionShell.scala 938:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"N/A"); // @[DandelionShell.scala 942:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_19) begin
          $fwrite(32'h80000002,"\n"); // @[DandelionShell.scala 944:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
