module LockingRRArbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [21:0] io_in_0_bits_address,
  input  [31:0] io_in_0_bits_data,
  input  [9:0]  io_in_0_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [21:0] io_out_bits_address,
  output [31:0] io_out_bits_data,
  output [9:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ,
  output        io_chosen
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? 1'h0 : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_address = io_chosen ? 22'h0 : io_in_0_bits_address; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? 32'h0 : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? 10'h0 : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_Typ = io_chosen ? 8'h0 : 8'h3; // @[Arbiter.scala 42:15]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 40:13]
endmodule
module ArbiterTree(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [21:0] io_in_0_bits_address,
  input  [31:0] io_in_0_bits_data,
  input  [9:0]  io_in_0_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [21:0] io_out_bits_address,
  output [31:0] io_out_bits_data,
  output [9:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ
);
  wire  LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_chosen; // @[ArbiterTree.scala 32:13]
  LockingRRArbiter LockingRRArbiter ( // @[ArbiterTree.scala 32:13]
    .io_in_0_ready(LockingRRArbiter_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_io_in_0_valid),
    .io_in_0_bits_address(LockingRRArbiter_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_io_in_0_bits_taskID),
    .io_out_ready(LockingRRArbiter_io_out_ready),
    .io_out_valid(LockingRRArbiter_io_out_valid),
    .io_out_bits_address(LockingRRArbiter_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_io_chosen)
  );
  assign io_in_0_ready = LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_out_valid = LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_address = LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_data = LockingRRArbiter_io_out_bits_data; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_taskID = LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_Typ = LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 65:12]
  assign LockingRRArbiter_io_in_0_valid = io_in_0_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_address = io_in_0_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_data = io_in_0_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_taskID = io_in_0_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_out_ready = io_out_ready; // @[ArbiterTree.scala 65:12]
endmodule
module Arbiter(
  output  io_in_0_ready,
  input   io_in_0_valid,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_out_ready,
  output  io_out_valid
);
  wire  _T_70; // @[Arbiter.scala 31:78]
  wire  _T_74; // @[Arbiter.scala 135:19]
  assign _T_70 = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_74 = _T_70 == 1'h0; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = _T_70 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_74 | io_in_1_valid; // @[Arbiter.scala 135:16]
endmodule
module Arbiter_1(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_data,
  input  [3:0]  io_in_0_bits_mask,
  input  [7:0]  io_in_0_bits_tag,
  input  [9:0]  io_in_0_bits_taskID,
  input         io_in_0_bits_iswrite,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_data,
  input  [3:0]  io_in_1_bits_mask,
  input  [7:0]  io_in_1_bits_tag,
  input  [9:0]  io_in_1_bits_taskID,
  input         io_in_1_bits_iswrite,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_data,
  output [3:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [9:0]  io_out_bits_taskID,
  output        io_out_bits_iswrite
);
  wire  _T_70; // @[Arbiter.scala 31:78]
  wire  _T_74; // @[Arbiter.scala 135:19]
  assign _T_70 = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_74 = _T_70 == 1'h0; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = _T_70 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_74 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_mask = io_in_0_valid ? io_in_0_bits_mask : io_in_1_bits_mask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_tag = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_taskID = io_in_0_valid ? io_in_0_bits_taskID : io_in_1_bits_taskID; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_iswrite = io_in_0_valid ? io_in_0_bits_iswrite : io_in_1_bits_iswrite; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Demux(
  input         io_en,
  input  [31:0] io_input_data,
  input  [7:0]  io_input_tag,
  input         io_sel,
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output [7:0]  io_outputs_0_tag,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data,
  output [7:0]  io_outputs_1_tag
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en ? _GEN_0 : 1'h0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_0_tag = io_input_tag; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en ? io_sel : 1'h0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_1_tag = io_input_tag; // @[Muxes.scala 23:19]
endmodule
module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output        io_chosen
);
  reg  _T_81; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  wire  _T_84; // @[Arbiter.scala 67:57]
  wire  _T_86; // @[Arbiter.scala 68:83]
  wire  _T_89; // @[Arbiter.scala 31:68]
  wire  _T_95; // @[Arbiter.scala 31:78]
  wire  _GEN_11; // @[Arbiter.scala 77:27]
  assign _T_84 = 1'h1 > _T_81; // @[Arbiter.scala 67:57]
  assign _T_86 = io_in_1_valid & _T_84; // @[Arbiter.scala 68:83]
  assign _T_89 = _T_86 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_95 = _T_89 == 1'h0; // @[Arbiter.scala 31:78]
  assign _GEN_11 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_86 == 1'h0; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_84 | _T_95; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_86 ? 1'h1 : _GEN_11; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_81 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_out_valid) begin
      _T_81 <= io_chosen;
    end
  end
endmodule
module Demux_1(
  input   io_en,
  input   io_sel,
  output  io_outputs_0_valid
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en ? _GEN_0 : 1'h0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
endmodule
module DeMuxTree(
  output        io_outputs_0_valid,
  input  [15:0] io_input_RouteID,
  input         io_enable
);
  wire  Demux_io_en; // @[Muxes.scala 91:13]
  wire  Demux_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_0_valid; // @[Muxes.scala 91:13]
  Demux_1 Demux ( // @[Muxes.scala 91:13]
    .io_en(Demux_io_en),
    .io_sel(Demux_io_sel),
    .io_outputs_0_valid(Demux_io_outputs_0_valid)
  );
  assign io_outputs_0_valid = Demux_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign Demux_io_en = io_enable; // @[Muxes.scala 135:14]
  assign Demux_io_sel = io_input_RouteID[0]; // @[Muxes.scala 136:15]
endmodule
module WriteTableEntry(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [21:0] io_NodeReq_bits_address,
  input  [31:0] io_NodeReq_bits_data,
  input  [9:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output        io_free
);
  reg [15:0] request_R_RouteID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_0;
  reg [9:0] request_R_taskID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_1;
  reg [7:0] sendbytemask; // @[WriteMemoryController.scala 61:29]
  reg [31:0] _RAND_2;
  reg [31:0] ReqAddress; // @[WriteMemoryController.scala 65:27]
  reg [31:0] _RAND_3;
  reg  ptr; // @[WriteMemoryController.scala 70:27]
  reg [31:0] _RAND_4;
  reg [31:0] linebuffer_0; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_5;
  reg [31:0] linebuffer_1; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_6;
  reg [1:0] state; // @[WriteMemoryController.scala 76:68]
  reg [31:0] _RAND_7;
  wire  _T_100; // @[WriteMemoryController.scala 89:21]
  wire [2:0] _T_106; // @[Cat.scala 30:58]
  wire [31:0] _GEN_29; // @[WriteMemoryController.scala 100:37]
  wire [32:0] _T_107; // @[WriteMemoryController.scala 100:37]
  reg  isWrite; // @[WriteMemoryController.scala 108:24]
  reg [31:0] _RAND_8;
  wire  _T_119; // @[Decoupled.scala 37:37]
  wire [19:0] _T_120; // @[WriteMemoryController.scala 121:44]
  wire [21:0] _GEN_30; // @[WriteMemoryController.scala 121:69]
  wire [21:0] _T_121; // @[WriteMemoryController.scala 121:69]
  wire  _T_122; // @[helpers.scala 27:24]
  wire  _T_123; // @[helpers.scala 27:47]
  wire  _T_124; // @[helpers.scala 27:40]
  wire  _T_130; // @[helpers.scala 28:15]
  wire  _T_131; // @[helpers.scala 28:38]
  wire  _T_132; // @[helpers.scala 28:31]
  wire  _T_138; // @[helpers.scala 29:17]
  wire  _T_139; // @[helpers.scala 29:40]
  wire  _T_140; // @[helpers.scala 29:33]
  wire [1:0] _T_154; // @[helpers.scala 39:32]
  wire [4:0] _T_156; // @[Cat.scala 30:58]
  wire [7:0] _T_183; // @[helpers.scala 50:12]
  wire [7:0] _T_184; // @[helpers.scala 49:10]
  wire [7:0] _T_185; // @[helpers.scala 48:19]
  wire [10:0] _GEN_32; // @[helpers.scala 20:26]
  wire [10:0] _T_187; // @[helpers.scala 20:26]
  wire [62:0] _GEN_33; // @[WriteMemoryController.scala 127:41]
  wire [62:0] _T_191; // @[WriteMemoryController.scala 127:41]
  wire [63:0] _T_209;
  wire [31:0] _T_210; // @[WriteMemoryController.scala 127:121]
  wire [31:0] _T_211; // @[WriteMemoryController.scala 127:121]
  wire [9:0] _GEN_3; // @[WriteMemoryController.scala 117:28]
  wire [15:0] _GEN_7; // @[WriteMemoryController.scala 117:28]
  wire [31:0] _GEN_8; // @[WriteMemoryController.scala 117:28]
  wire [10:0] _GEN_10; // @[WriteMemoryController.scala 117:28]
  wire [31:0] _GEN_11; // @[WriteMemoryController.scala 117:28]
  wire [31:0] _GEN_12; // @[WriteMemoryController.scala 117:28]
  wire [1:0] _GEN_13; // @[WriteMemoryController.scala 117:28]
  wire  _T_212; // @[WriteMemoryController.scala 139:15]
  wire  _T_214; // @[WriteMemoryController.scala 139:47]
  wire  _T_215; // @[WriteMemoryController.scala 139:30]
  wire  _T_217; // @[Decoupled.scala 37:37]
  wire [3:0] _T_218; // @[WriteMemoryController.scala 144:36]
  wire [1:0] _T_220; // @[WriteMemoryController.scala 146:18]
  wire  _T_221; // @[WriteMemoryController.scala 146:18]
  wire [10:0] _GEN_14; // @[WriteMemoryController.scala 142:29]
  wire  _GEN_15; // @[WriteMemoryController.scala 142:29]
  wire [1:0] _GEN_16; // @[WriteMemoryController.scala 142:29]
  wire [10:0] _GEN_18; // @[WriteMemoryController.scala 139:76]
  wire  _GEN_19; // @[WriteMemoryController.scala 139:76]
  wire [1:0] _GEN_20; // @[WriteMemoryController.scala 139:76]
  wire  _T_222; // @[WriteMemoryController.scala 156:15]
  wire  _T_225; // @[WriteMemoryController.scala 156:32]
  wire  _T_227; // @[WriteMemoryController.scala 158:27]
  wire [1:0] _T_228; // @[WriteMemoryController.scala 159:17]
  wire [1:0] _GEN_21; // @[WriteMemoryController.scala 156:66]
  wire  _T_233; // @[Decoupled.scala 37:37]
  wire [1:0] _GEN_22; // @[WriteMemoryController.scala 173:29]
  wire  _GEN_25; // @[WriteMemoryController.scala 166:26]
  wire [1:0] _GEN_27; // @[WriteMemoryController.scala 166:26]
  assign _T_100 = state == 2'h3; // @[WriteMemoryController.scala 89:21]
  assign _T_106 = {ptr,2'h0}; // @[Cat.scala 30:58]
  assign _GEN_29 = {{29'd0}, _T_106}; // @[WriteMemoryController.scala 100:37]
  assign _T_107 = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:37]
  assign _T_119 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 37:37]
  assign _T_120 = io_NodeReq_bits_address[21:2]; // @[WriteMemoryController.scala 121:44]
  assign _GEN_30 = {{2'd0}, _T_120}; // @[WriteMemoryController.scala 121:69]
  assign _T_121 = _GEN_30 << 2; // @[WriteMemoryController.scala 121:69]
  assign _T_122 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_123 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_124 = _T_122 | _T_123; // @[helpers.scala 27:40]
  assign _T_130 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_131 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_132 = _T_130 | _T_131; // @[helpers.scala 28:31]
  assign _T_138 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_139 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_140 = _T_138 | _T_139; // @[helpers.scala 29:33]
  assign _T_154 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_156 = {_T_154,3'h0}; // @[Cat.scala 30:58]
  assign _T_183 = _T_140 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_184 = _T_132 ? 8'h1 : _T_183; // @[helpers.scala 49:10]
  assign _T_185 = _T_124 ? 8'h3 : _T_184; // @[helpers.scala 48:19]
  assign _GEN_32 = {{3'd0}, _T_185}; // @[helpers.scala 20:26]
  assign _T_187 = _GEN_32 << _T_154; // @[helpers.scala 20:26]
  assign _GEN_33 = {{31'd0}, io_NodeReq_bits_data}; // @[WriteMemoryController.scala 127:41]
  assign _T_191 = _GEN_33 << _T_156; // @[WriteMemoryController.scala 127:41]
  assign _T_209 = {{1'd0}, _T_191};
  assign _T_210 = _T_209[31:0]; // @[WriteMemoryController.scala 127:121]
  assign _T_211 = _T_209[63:32]; // @[WriteMemoryController.scala 127:121]
  assign _GEN_3 = _T_119 ? io_NodeReq_bits_taskID : request_R_taskID; // @[WriteMemoryController.scala 117:28]
  assign _GEN_7 = _T_119 ? 16'h0 : request_R_RouteID; // @[WriteMemoryController.scala 117:28]
  assign _GEN_8 = _T_119 ? {{10'd0}, _T_121} : ReqAddress; // @[WriteMemoryController.scala 117:28]
  assign _GEN_10 = _T_119 ? _T_187 : {{3'd0}, sendbytemask}; // @[WriteMemoryController.scala 117:28]
  assign _GEN_11 = _T_119 ? _T_210 : linebuffer_0; // @[WriteMemoryController.scala 117:28]
  assign _GEN_12 = _T_119 ? _T_211 : linebuffer_1; // @[WriteMemoryController.scala 117:28]
  assign _GEN_13 = _T_119 ? 2'h1 : state; // @[WriteMemoryController.scala 117:28]
  assign _T_212 = state == 2'h1; // @[WriteMemoryController.scala 139:15]
  assign _T_214 = sendbytemask != 8'h0; // @[WriteMemoryController.scala 139:47]
  assign _T_215 = _T_212 & _T_214; // @[WriteMemoryController.scala 139:30]
  assign _T_217 = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 37:37]
  assign _T_218 = sendbytemask[7:4]; // @[WriteMemoryController.scala 144:36]
  assign _T_220 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _T_221 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _GEN_14 = _T_217 ? {{7'd0}, _T_218} : _GEN_10; // @[WriteMemoryController.scala 142:29]
  assign _GEN_15 = _T_217 ? _T_221 : ptr; // @[WriteMemoryController.scala 142:29]
  assign _GEN_16 = _T_217 ? 2'h2 : _GEN_13; // @[WriteMemoryController.scala 142:29]
  assign _GEN_18 = _T_215 ? _GEN_14 : _GEN_10; // @[WriteMemoryController.scala 139:76]
  assign _GEN_19 = _T_215 ? _GEN_15 : ptr; // @[WriteMemoryController.scala 139:76]
  assign _GEN_20 = _T_215 ? _GEN_16 : _GEN_13; // @[WriteMemoryController.scala 139:76]
  assign _T_222 = state == 2'h2; // @[WriteMemoryController.scala 156:15]
  assign _T_225 = _T_222 & io_MemResp_valid; // @[WriteMemoryController.scala 156:32]
  assign _T_227 = sendbytemask == 8'h0; // @[WriteMemoryController.scala 158:27]
  assign _T_228 = _T_227 ? 2'h3 : 2'h1; // @[WriteMemoryController.scala 159:17]
  assign _GEN_21 = _T_225 ? _T_228 : _GEN_20; // @[WriteMemoryController.scala 156:66]
  assign _T_233 = io_output_ready & io_output_valid; // @[Decoupled.scala 37:37]
  assign _GEN_22 = _T_233 ? 2'h0 : _GEN_21; // @[WriteMemoryController.scala 173:29]
  assign _GEN_25 = _T_100 ? 1'h0 : _GEN_19; // @[WriteMemoryController.scala 166:26]
  assign _GEN_27 = _T_100 ? _GEN_22 : _GEN_21; // @[WriteMemoryController.scala 166:26]
  assign io_NodeReq_ready = state == 2'h0; // @[WriteMemoryController.scala 87:20]
  assign io_MemReq_valid = _T_212 & _T_214; // @[WriteMemoryController.scala 99:19 WriteMemoryController.scala 140:21]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:23]
  assign io_MemReq_bits_data = ptr ? linebuffer_1 : linebuffer_0; // @[WriteMemoryController.scala 102:23]
  assign io_MemReq_bits_mask = sendbytemask[3:0]; // @[WriteMemoryController.scala 103:23]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[WriteMemoryController.scala 110:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[WriteMemoryController.scala 109:26]
  assign io_output_valid = state == 2'h3; // @[WriteMemoryController.scala 95:19 WriteMemoryController.scala 168:21]
  assign io_output_bits_RouteID = request_R_RouteID; // @[WriteMemoryController.scala 98:26]
  assign io_free = state == 2'h0; // @[WriteMemoryController.scala 85:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  request_R_RouteID = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_taskID = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sendbytemask = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ReqAddress = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ptr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  linebuffer_0 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  linebuffer_1 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  isWrite = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_119) begin
        request_R_RouteID <= 16'h0;
      end
    end
    if (reset) begin
      request_R_taskID <= 10'h0;
    end else begin
      if (_T_119) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_18[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_119) begin
        ReqAddress <= {{10'd0}, _T_121};
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (_T_100) begin
        ptr <= 1'h0;
      end else begin
        if (_T_215) begin
          if (_T_217) begin
            ptr <= _T_221;
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (_T_119) begin
        linebuffer_0 <= _T_210;
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (_T_119) begin
        linebuffer_1 <= _T_211;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_100) begin
        if (_T_233) begin
          state <= 2'h0;
        end else begin
          if (_T_225) begin
            if (_T_227) begin
              state <= 2'h3;
            end else begin
              state <= 2'h1;
            end
          end else begin
            if (_T_215) begin
              if (_T_217) begin
                state <= 2'h2;
              end else begin
                if (_T_119) begin
                  state <= 2'h1;
                end
              end
            end else begin
              if (_T_119) begin
                state <= 2'h1;
              end
            end
          end
        end
      end else begin
        if (_T_225) begin
          if (_T_227) begin
            state <= 2'h3;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_215) begin
            if (_T_217) begin
              state <= 2'h2;
            end else begin
              if (_T_119) begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_119) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      isWrite <= 1'h0;
    end else begin
      isWrite <= 1'h1;
    end
  end
endmodule
module WriteTableEntry_1(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [21:0] io_NodeReq_bits_address,
  input  [31:0] io_NodeReq_bits_data,
  input  [9:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output        io_free
);
  reg [15:0] request_R_RouteID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_0;
  reg [9:0] request_R_taskID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_1;
  reg [7:0] sendbytemask; // @[WriteMemoryController.scala 61:29]
  reg [31:0] _RAND_2;
  reg [31:0] ReqAddress; // @[WriteMemoryController.scala 65:27]
  reg [31:0] _RAND_3;
  reg  ptr; // @[WriteMemoryController.scala 70:27]
  reg [31:0] _RAND_4;
  reg [31:0] linebuffer_0; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_5;
  reg [31:0] linebuffer_1; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_6;
  reg [1:0] state; // @[WriteMemoryController.scala 76:68]
  reg [31:0] _RAND_7;
  wire  _T_92; // @[WriteMemoryController.scala 89:21]
  wire [2:0] _T_98; // @[Cat.scala 30:58]
  wire [31:0] _GEN_29; // @[WriteMemoryController.scala 100:37]
  wire [32:0] _T_99; // @[WriteMemoryController.scala 100:37]
  reg  myID; // @[WriteMemoryController.scala 106:21]
  reg [31:0] _RAND_8;
  reg  isWrite; // @[WriteMemoryController.scala 108:24]
  reg [31:0] _RAND_9;
  wire  _T_111; // @[Decoupled.scala 37:37]
  wire [19:0] _T_112; // @[WriteMemoryController.scala 121:44]
  wire [21:0] _GEN_30; // @[WriteMemoryController.scala 121:69]
  wire [21:0] _T_113; // @[WriteMemoryController.scala 121:69]
  wire  _T_114; // @[helpers.scala 27:24]
  wire  _T_115; // @[helpers.scala 27:47]
  wire  _T_116; // @[helpers.scala 27:40]
  wire  _T_122; // @[helpers.scala 28:15]
  wire  _T_123; // @[helpers.scala 28:38]
  wire  _T_124; // @[helpers.scala 28:31]
  wire  _T_130; // @[helpers.scala 29:17]
  wire  _T_131; // @[helpers.scala 29:40]
  wire  _T_132; // @[helpers.scala 29:33]
  wire [1:0] _T_146; // @[helpers.scala 39:32]
  wire [4:0] _T_148; // @[Cat.scala 30:58]
  wire [7:0] _T_175; // @[helpers.scala 50:12]
  wire [7:0] _T_176; // @[helpers.scala 49:10]
  wire [7:0] _T_177; // @[helpers.scala 48:19]
  wire [10:0] _GEN_32; // @[helpers.scala 20:26]
  wire [10:0] _T_179; // @[helpers.scala 20:26]
  wire [62:0] _GEN_33; // @[WriteMemoryController.scala 127:41]
  wire [62:0] _T_183; // @[WriteMemoryController.scala 127:41]
  wire [63:0] _T_201;
  wire [31:0] _T_202; // @[WriteMemoryController.scala 127:121]
  wire [31:0] _T_203; // @[WriteMemoryController.scala 127:121]
  wire [9:0] _GEN_3; // @[WriteMemoryController.scala 117:28]
  wire [15:0] _GEN_7; // @[WriteMemoryController.scala 117:28]
  wire [31:0] _GEN_8; // @[WriteMemoryController.scala 117:28]
  wire [10:0] _GEN_10; // @[WriteMemoryController.scala 117:28]
  wire [31:0] _GEN_11; // @[WriteMemoryController.scala 117:28]
  wire [31:0] _GEN_12; // @[WriteMemoryController.scala 117:28]
  wire [1:0] _GEN_13; // @[WriteMemoryController.scala 117:28]
  wire  _T_204; // @[WriteMemoryController.scala 139:15]
  wire  _T_206; // @[WriteMemoryController.scala 139:47]
  wire  _T_207; // @[WriteMemoryController.scala 139:30]
  wire  _T_209; // @[Decoupled.scala 37:37]
  wire [3:0] _T_210; // @[WriteMemoryController.scala 144:36]
  wire [1:0] _T_212; // @[WriteMemoryController.scala 146:18]
  wire  _T_213; // @[WriteMemoryController.scala 146:18]
  wire [10:0] _GEN_14; // @[WriteMemoryController.scala 142:29]
  wire  _GEN_15; // @[WriteMemoryController.scala 142:29]
  wire [1:0] _GEN_16; // @[WriteMemoryController.scala 142:29]
  wire [10:0] _GEN_18; // @[WriteMemoryController.scala 139:76]
  wire  _GEN_19; // @[WriteMemoryController.scala 139:76]
  wire [1:0] _GEN_20; // @[WriteMemoryController.scala 139:76]
  wire  _T_214; // @[WriteMemoryController.scala 156:15]
  wire  _T_217; // @[WriteMemoryController.scala 156:32]
  wire  _T_219; // @[WriteMemoryController.scala 158:27]
  wire [1:0] _T_220; // @[WriteMemoryController.scala 159:17]
  wire [1:0] _GEN_21; // @[WriteMemoryController.scala 156:66]
  wire  _T_225; // @[Decoupled.scala 37:37]
  wire [1:0] _GEN_22; // @[WriteMemoryController.scala 173:29]
  wire  _GEN_25; // @[WriteMemoryController.scala 166:26]
  wire [1:0] _GEN_27; // @[WriteMemoryController.scala 166:26]
  assign _T_92 = state == 2'h3; // @[WriteMemoryController.scala 89:21]
  assign _T_98 = {ptr,2'h0}; // @[Cat.scala 30:58]
  assign _GEN_29 = {{29'd0}, _T_98}; // @[WriteMemoryController.scala 100:37]
  assign _T_99 = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:37]
  assign _T_111 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 37:37]
  assign _T_112 = io_NodeReq_bits_address[21:2]; // @[WriteMemoryController.scala 121:44]
  assign _GEN_30 = {{2'd0}, _T_112}; // @[WriteMemoryController.scala 121:69]
  assign _T_113 = _GEN_30 << 2; // @[WriteMemoryController.scala 121:69]
  assign _T_114 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_115 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_116 = _T_114 | _T_115; // @[helpers.scala 27:40]
  assign _T_122 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_123 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_124 = _T_122 | _T_123; // @[helpers.scala 28:31]
  assign _T_130 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_131 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_132 = _T_130 | _T_131; // @[helpers.scala 29:33]
  assign _T_146 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_148 = {_T_146,3'h0}; // @[Cat.scala 30:58]
  assign _T_175 = _T_132 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_176 = _T_124 ? 8'h1 : _T_175; // @[helpers.scala 49:10]
  assign _T_177 = _T_116 ? 8'h3 : _T_176; // @[helpers.scala 48:19]
  assign _GEN_32 = {{3'd0}, _T_177}; // @[helpers.scala 20:26]
  assign _T_179 = _GEN_32 << _T_146; // @[helpers.scala 20:26]
  assign _GEN_33 = {{31'd0}, io_NodeReq_bits_data}; // @[WriteMemoryController.scala 127:41]
  assign _T_183 = _GEN_33 << _T_148; // @[WriteMemoryController.scala 127:41]
  assign _T_201 = {{1'd0}, _T_183};
  assign _T_202 = _T_201[31:0]; // @[WriteMemoryController.scala 127:121]
  assign _T_203 = _T_201[63:32]; // @[WriteMemoryController.scala 127:121]
  assign _GEN_3 = _T_111 ? io_NodeReq_bits_taskID : request_R_taskID; // @[WriteMemoryController.scala 117:28]
  assign _GEN_7 = _T_111 ? 16'h0 : request_R_RouteID; // @[WriteMemoryController.scala 117:28]
  assign _GEN_8 = _T_111 ? {{10'd0}, _T_113} : ReqAddress; // @[WriteMemoryController.scala 117:28]
  assign _GEN_10 = _T_111 ? _T_179 : {{3'd0}, sendbytemask}; // @[WriteMemoryController.scala 117:28]
  assign _GEN_11 = _T_111 ? _T_202 : linebuffer_0; // @[WriteMemoryController.scala 117:28]
  assign _GEN_12 = _T_111 ? _T_203 : linebuffer_1; // @[WriteMemoryController.scala 117:28]
  assign _GEN_13 = _T_111 ? 2'h1 : state; // @[WriteMemoryController.scala 117:28]
  assign _T_204 = state == 2'h1; // @[WriteMemoryController.scala 139:15]
  assign _T_206 = sendbytemask != 8'h0; // @[WriteMemoryController.scala 139:47]
  assign _T_207 = _T_204 & _T_206; // @[WriteMemoryController.scala 139:30]
  assign _T_209 = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 37:37]
  assign _T_210 = sendbytemask[7:4]; // @[WriteMemoryController.scala 144:36]
  assign _T_212 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _T_213 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _GEN_14 = _T_209 ? {{7'd0}, _T_210} : _GEN_10; // @[WriteMemoryController.scala 142:29]
  assign _GEN_15 = _T_209 ? _T_213 : ptr; // @[WriteMemoryController.scala 142:29]
  assign _GEN_16 = _T_209 ? 2'h2 : _GEN_13; // @[WriteMemoryController.scala 142:29]
  assign _GEN_18 = _T_207 ? _GEN_14 : _GEN_10; // @[WriteMemoryController.scala 139:76]
  assign _GEN_19 = _T_207 ? _GEN_15 : ptr; // @[WriteMemoryController.scala 139:76]
  assign _GEN_20 = _T_207 ? _GEN_16 : _GEN_13; // @[WriteMemoryController.scala 139:76]
  assign _T_214 = state == 2'h2; // @[WriteMemoryController.scala 156:15]
  assign _T_217 = _T_214 & io_MemResp_valid; // @[WriteMemoryController.scala 156:32]
  assign _T_219 = sendbytemask == 8'h0; // @[WriteMemoryController.scala 158:27]
  assign _T_220 = _T_219 ? 2'h3 : 2'h1; // @[WriteMemoryController.scala 159:17]
  assign _GEN_21 = _T_217 ? _T_220 : _GEN_20; // @[WriteMemoryController.scala 156:66]
  assign _T_225 = io_output_ready & io_output_valid; // @[Decoupled.scala 37:37]
  assign _GEN_22 = _T_225 ? 2'h0 : _GEN_21; // @[WriteMemoryController.scala 173:29]
  assign _GEN_25 = _T_92 ? 1'h0 : _GEN_19; // @[WriteMemoryController.scala 166:26]
  assign _GEN_27 = _T_92 ? _GEN_22 : _GEN_21; // @[WriteMemoryController.scala 166:26]
  assign io_NodeReq_ready = state == 2'h0; // @[WriteMemoryController.scala 87:20]
  assign io_MemReq_valid = _T_204 & _T_206; // @[WriteMemoryController.scala 99:19 WriteMemoryController.scala 140:21]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:23]
  assign io_MemReq_bits_data = ptr ? linebuffer_1 : linebuffer_0; // @[WriteMemoryController.scala 102:23]
  assign io_MemReq_bits_mask = sendbytemask[3:0]; // @[WriteMemoryController.scala 103:23]
  assign io_MemReq_bits_tag = {{7'd0}, myID}; // @[WriteMemoryController.scala 107:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[WriteMemoryController.scala 110:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[WriteMemoryController.scala 109:26]
  assign io_output_valid = state == 2'h3; // @[WriteMemoryController.scala 95:19 WriteMemoryController.scala 168:21]
  assign io_output_bits_RouteID = request_R_RouteID; // @[WriteMemoryController.scala 98:26]
  assign io_free = state == 2'h0; // @[WriteMemoryController.scala 85:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  request_R_RouteID = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_taskID = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sendbytemask = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ReqAddress = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ptr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  linebuffer_0 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  linebuffer_1 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  myID = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  isWrite = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_111) begin
        request_R_RouteID <= 16'h0;
      end
    end
    if (reset) begin
      request_R_taskID <= 10'h0;
    end else begin
      if (_T_111) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_18[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_111) begin
        ReqAddress <= {{10'd0}, _T_113};
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (_T_92) begin
        ptr <= 1'h0;
      end else begin
        if (_T_207) begin
          if (_T_209) begin
            ptr <= _T_213;
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (_T_111) begin
        linebuffer_0 <= _T_202;
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (_T_111) begin
        linebuffer_1 <= _T_203;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_92) begin
        if (_T_225) begin
          state <= 2'h0;
        end else begin
          if (_T_217) begin
            if (_T_219) begin
              state <= 2'h3;
            end else begin
              state <= 2'h1;
            end
          end else begin
            if (_T_207) begin
              if (_T_209) begin
                state <= 2'h2;
              end else begin
                if (_T_111) begin
                  state <= 2'h1;
                end
              end
            end else begin
              if (_T_111) begin
                state <= 2'h1;
              end
            end
          end
        end
      end else begin
        if (_T_217) begin
          if (_T_219) begin
            state <= 2'h3;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_207) begin
            if (_T_209) begin
              state <= 2'h2;
            end else begin
              if (_T_111) begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_111) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      myID <= 1'h0;
    end else begin
      myID <= 1'h1;
    end
    if (reset) begin
      isWrite <= 1'h0;
    end else begin
      isWrite <= 1'h1;
    end
  end
endmodule
module WriteMemoryController(
  input         clock,
  input         reset,
  output        io_WriteIn_0_ready,
  input         io_WriteIn_0_valid,
  input  [21:0] io_WriteIn_0_bits_address,
  input  [31:0] io_WriteIn_0_bits_data,
  input  [9:0]  io_WriteIn_0_bits_taskID,
  output        io_WriteOut_0_valid,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag
);
  wire  in_arb_io_in_0_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_0_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_0_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_0_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [9:0] in_arb_io_in_0_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_out_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_out_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_out_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_out_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [9:0] in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire [7:0] in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 194:25]
  wire  alloc_arb_io_in_0_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_0_valid; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_1_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_1_valid; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_out_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_out_valid; // @[WriteMemoryController.scala 196:25]
  wire  cachereq_arb_io_in_0_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_0_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [9:0] cachereq_arb_io_in_0_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [9:0] cachereq_arb_io_in_1_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [9:0] cachereq_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cacheresp_demux_io_en; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_sel; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[WriteMemoryController.scala 201:31]
  wire  out_arb_clock; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_0_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_0_valid; // @[WriteMemoryController.scala 204:25]
  wire [15:0] out_arb_io_in_0_bits_RouteID; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_1_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_1_valid; // @[WriteMemoryController.scala 204:25]
  wire [15:0] out_arb_io_in_1_bits_RouteID; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_out_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_out_valid; // @[WriteMemoryController.scala 204:25]
  wire [15:0] out_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_chosen; // @[WriteMemoryController.scala 204:25]
  wire  out_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 205:25]
  wire [15:0] out_demux_io_input_RouteID; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_enable; // @[WriteMemoryController.scala 205:25]
  wire  WriteTable_0_clock; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_reset; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_NodeReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_NodeReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [21:0] WriteTable_0_io_NodeReq_bits_address; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_NodeReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [9:0] WriteTable_0_io_NodeReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_0_io_NodeReq_bits_Typ; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_MemReq_bits_addr; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_MemReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [3:0] WriteTable_0_io_MemReq_bits_mask; // @[WriteMemoryController.scala 223:29]
  wire [9:0] WriteTable_0_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemResp_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_output_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_output_valid; // @[WriteMemoryController.scala 223:29]
  wire [15:0] WriteTable_0_io_output_bits_RouteID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_free; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_clock; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_reset; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_NodeReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_NodeReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [21:0] WriteTable_1_io_NodeReq_bits_address; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_NodeReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [9:0] WriteTable_1_io_NodeReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_1_io_NodeReq_bits_Typ; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_MemReq_bits_addr; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_MemReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [3:0] WriteTable_1_io_MemReq_bits_mask; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_1_io_MemReq_bits_tag; // @[WriteMemoryController.scala 223:29]
  wire [9:0] WriteTable_1_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemResp_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_output_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_output_valid; // @[WriteMemoryController.scala 223:29]
  wire [15:0] WriteTable_1_io_output_bits_RouteID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_free; // @[WriteMemoryController.scala 223:29]
  ArbiterTree in_arb ( // @[WriteMemoryController.scala 194:25]
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_address(in_arb_io_in_0_bits_address),
    .io_in_0_bits_data(in_arb_io_in_0_bits_data),
    .io_in_0_bits_taskID(in_arb_io_in_0_bits_taskID),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_address(in_arb_io_out_bits_address),
    .io_out_bits_data(in_arb_io_out_bits_data),
    .io_out_bits_taskID(in_arb_io_out_bits_taskID),
    .io_out_bits_Typ(in_arb_io_out_bits_Typ)
  );
  Arbiter alloc_arb ( // @[WriteMemoryController.scala 196:25]
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid)
  );
  Arbiter_1 cachereq_arb ( // @[WriteMemoryController.scala 199:31]
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite)
  );
  Demux cacheresp_demux ( // @[WriteMemoryController.scala 201:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  RRArbiter out_arb ( // @[WriteMemoryController.scala 204:25]
    .clock(out_arb_clock),
    .io_in_0_ready(out_arb_io_in_0_ready),
    .io_in_0_valid(out_arb_io_in_0_valid),
    .io_in_0_bits_RouteID(out_arb_io_in_0_bits_RouteID),
    .io_in_1_ready(out_arb_io_in_1_ready),
    .io_in_1_valid(out_arb_io_in_1_valid),
    .io_in_1_bits_RouteID(out_arb_io_in_1_bits_RouteID),
    .io_out_ready(out_arb_io_out_ready),
    .io_out_valid(out_arb_io_out_valid),
    .io_out_bits_RouteID(out_arb_io_out_bits_RouteID),
    .io_chosen(out_arb_io_chosen)
  );
  DeMuxTree out_demux ( // @[WriteMemoryController.scala 205:25]
    .io_outputs_0_valid(out_demux_io_outputs_0_valid),
    .io_input_RouteID(out_demux_io_input_RouteID),
    .io_enable(out_demux_io_enable)
  );
  WriteTableEntry WriteTable_0 ( // @[WriteMemoryController.scala 223:29]
    .clock(WriteTable_0_clock),
    .reset(WriteTable_0_reset),
    .io_NodeReq_ready(WriteTable_0_io_NodeReq_ready),
    .io_NodeReq_valid(WriteTable_0_io_NodeReq_valid),
    .io_NodeReq_bits_address(WriteTable_0_io_NodeReq_bits_address),
    .io_NodeReq_bits_data(WriteTable_0_io_NodeReq_bits_data),
    .io_NodeReq_bits_taskID(WriteTable_0_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(WriteTable_0_io_NodeReq_bits_Typ),
    .io_MemReq_ready(WriteTable_0_io_MemReq_ready),
    .io_MemReq_valid(WriteTable_0_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteTable_0_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteTable_0_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteTable_0_io_MemReq_bits_mask),
    .io_MemReq_bits_taskID(WriteTable_0_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteTable_0_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteTable_0_io_MemResp_valid),
    .io_output_ready(WriteTable_0_io_output_ready),
    .io_output_valid(WriteTable_0_io_output_valid),
    .io_output_bits_RouteID(WriteTable_0_io_output_bits_RouteID),
    .io_free(WriteTable_0_io_free)
  );
  WriteTableEntry_1 WriteTable_1 ( // @[WriteMemoryController.scala 223:29]
    .clock(WriteTable_1_clock),
    .reset(WriteTable_1_reset),
    .io_NodeReq_ready(WriteTable_1_io_NodeReq_ready),
    .io_NodeReq_valid(WriteTable_1_io_NodeReq_valid),
    .io_NodeReq_bits_address(WriteTable_1_io_NodeReq_bits_address),
    .io_NodeReq_bits_data(WriteTable_1_io_NodeReq_bits_data),
    .io_NodeReq_bits_taskID(WriteTable_1_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(WriteTable_1_io_NodeReq_bits_Typ),
    .io_MemReq_ready(WriteTable_1_io_MemReq_ready),
    .io_MemReq_valid(WriteTable_1_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteTable_1_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteTable_1_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteTable_1_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(WriteTable_1_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(WriteTable_1_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteTable_1_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteTable_1_io_MemResp_valid),
    .io_output_ready(WriteTable_1_io_output_ready),
    .io_output_valid(WriteTable_1_io_output_valid),
    .io_output_bits_RouteID(WriteTable_1_io_output_bits_RouteID),
    .io_free(WriteTable_1_io_free)
  );
  assign io_WriteIn_0_ready = in_arb_io_in_0_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteOut_0_valid = out_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 214:20]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[WriteMemoryController.scala 261:13]
  assign in_arb_io_in_0_valid = io_WriteIn_0_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_address = io_WriteIn_0_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_data = io_WriteIn_0_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_taskID = io_WriteIn_0_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_out_ready = alloc_arb_io_out_valid; // @[WriteMemoryController.scala 256:23]
  assign alloc_arb_io_in_0_valid = WriteTable_0_io_free; // @[WriteMemoryController.scala 226:30]
  assign alloc_arb_io_in_1_valid = WriteTable_1_io_free; // @[WriteMemoryController.scala 226:30]
  assign alloc_arb_io_out_ready = in_arb_io_out_valid; // @[WriteMemoryController.scala 257:26]
  assign cachereq_arb_io_in_0_valid = WriteTable_0_io_MemReq_valid; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_addr = WriteTable_0_io_MemReq_bits_addr; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_data = WriteTable_0_io_MemReq_bits_data; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_mask = WriteTable_0_io_MemReq_bits_mask; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_tag = 8'h0; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_taskID = WriteTable_0_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_iswrite = WriteTable_0_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_valid = WriteTable_1_io_MemReq_valid; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_addr = WriteTable_1_io_MemReq_bits_addr; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_data = WriteTable_1_io_MemReq_bits_data; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_mask = WriteTable_1_io_MemReq_bits_mask; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_tag = WriteTable_1_io_MemReq_bits_tag; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_taskID = WriteTable_1_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_iswrite = WriteTable_1_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[WriteMemoryController.scala 261:13]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[WriteMemoryController.scala 264:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[WriteMemoryController.scala 265:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[WriteMemoryController.scala 265:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_tag[0]; // @[WriteMemoryController.scala 266:26]
  assign out_arb_clock = clock;
  assign out_arb_io_in_0_valid = WriteTable_0_io_output_valid; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_0_bits_RouteID = WriteTable_0_io_output_bits_RouteID; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_1_valid = WriteTable_1_io_output_valid; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_1_bits_RouteID = WriteTable_1_io_output_bits_RouteID; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_out_ready = 1'h1; // @[WriteMemoryController.scala 269:24]
  assign out_demux_io_input_RouteID = out_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 271:22]
  assign out_demux_io_enable = out_arb_io_out_ready & out_arb_io_out_valid; // @[WriteMemoryController.scala 270:23]
  assign WriteTable_0_clock = clock;
  assign WriteTable_0_reset = reset;
  assign WriteTable_0_io_NodeReq_valid = alloc_arb_io_in_0_ready & alloc_arb_io_in_0_valid; // @[WriteMemoryController.scala 228:34]
  assign WriteTable_0_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_data = in_arb_io_out_bits_data; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_MemReq_ready = cachereq_arb_io_in_0_ready; // @[WriteMemoryController.scala 232:27]
  assign WriteTable_0_io_MemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 235:28]
  assign WriteTable_0_io_output_ready = out_arb_io_in_0_ready; // @[WriteMemoryController.scala 238:22]
  assign WriteTable_1_clock = clock;
  assign WriteTable_1_reset = reset;
  assign WriteTable_1_io_NodeReq_valid = alloc_arb_io_in_1_ready & alloc_arb_io_in_1_valid; // @[WriteMemoryController.scala 228:34]
  assign WriteTable_1_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_data = in_arb_io_out_bits_data; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_MemReq_ready = cachereq_arb_io_in_1_ready; // @[WriteMemoryController.scala 232:27]
  assign WriteTable_1_io_MemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 235:28]
  assign WriteTable_1_io_output_ready = out_arb_io_in_1_ready; // @[WriteMemoryController.scala 238:22]
endmodule
module LockingRRArbiter_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  input  [31:0] io_in_0_bits_address,
  input  [9:0]  io_in_0_bits_taskID,
  input  [7:0]  io_in_0_bits_Typ,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input  [31:0] io_in_1_bits_address,
  input  [9:0]  io_in_1_bits_taskID,
  input  [7:0]  io_in_1_bits_Typ,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_address,
  output [9:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ,
  output        io_chosen
);
  wire  _T_79; // @[Decoupled.scala 37:37]
  reg  _T_81; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  wire  _T_84; // @[Arbiter.scala 67:57]
  wire  _T_86; // @[Arbiter.scala 68:83]
  wire  _T_89; // @[Arbiter.scala 31:68]
  wire  _T_93; // @[Arbiter.scala 31:78]
  wire  _T_95; // @[Arbiter.scala 31:78]
  wire  _T_99; // @[Arbiter.scala 72:50]
  wire  _GEN_13; // @[Arbiter.scala 77:27]
  assign _T_79 = io_out_ready & io_out_valid; // @[Decoupled.scala 37:37]
  assign _T_84 = 1'h1 > _T_81; // @[Arbiter.scala 67:57]
  assign _T_86 = io_in_1_valid & _T_84; // @[Arbiter.scala 68:83]
  assign _T_89 = _T_86 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_93 = _T_86 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_95 = _T_89 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_99 = _T_84 | _T_95; // @[Arbiter.scala 72:50]
  assign _GEN_13 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_93 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_99 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_out_bits_address = io_chosen ? io_in_1_bits_address : io_in_0_bits_address; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_Typ = io_chosen ? io_in_1_bits_Typ : io_in_0_bits_Typ; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_86 ? 1'h1 : _GEN_13; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_81 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_79) begin
      _T_81 <= io_chosen;
    end
  end
endmodule
module ArbiterTree_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_address,
  input  [9:0]  io_in_0_bits_taskID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_address,
  input  [9:0]  io_in_1_bits_taskID,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_address,
  input  [9:0]  io_in_2_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_address,
  output [9:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ
);
  wire  LockingRRArbiter_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_1_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_1_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_1_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_2_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_2_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [9:0] LockingRRArbiter_2_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_chosen; // @[ArbiterTree.scala 32:13]
  LockingRRArbiter_1 LockingRRArbiter ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_clock),
    .io_in_0_ready(LockingRRArbiter_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_io_out_ready),
    .io_out_valid(LockingRRArbiter_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_io_chosen)
  );
  LockingRRArbiter_1 LockingRRArbiter_1 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_1_clock),
    .io_in_0_ready(LockingRRArbiter_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_1_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_1_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_1_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_1_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_1_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_1_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_1_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_1_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_1_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_1_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_1_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_1_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_1_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_1_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_1_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_1_io_chosen)
  );
  LockingRRArbiter_1 LockingRRArbiter_2 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_2_clock),
    .io_in_0_ready(LockingRRArbiter_2_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_2_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_2_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_2_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_2_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_2_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_2_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_2_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_2_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_2_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_2_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_2_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_2_io_out_ready),
    .io_out_valid(LockingRRArbiter_2_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_2_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_2_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_2_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_2_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_2_io_chosen)
  );
  assign io_in_0_ready = LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_1_ready = LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_2_ready = LockingRRArbiter_1_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_out_valid = LockingRRArbiter_2_io_out_valid; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_RouteID = LockingRRArbiter_2_io_out_bits_RouteID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_address = LockingRRArbiter_2_io_out_bits_address; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_taskID = LockingRRArbiter_2_io_out_bits_taskID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_Typ = LockingRRArbiter_2_io_out_bits_Typ; // @[ArbiterTree.scala 65:12]
  assign LockingRRArbiter_clock = clock;
  assign LockingRRArbiter_io_in_0_valid = io_in_0_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_RouteID = 16'h0; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_address = io_in_0_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_taskID = io_in_0_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_valid = io_in_1_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_RouteID = 16'h1; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_address = io_in_1_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_taskID = io_in_1_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_out_ready = LockingRRArbiter_2_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_1_clock = clock;
  assign LockingRRArbiter_1_io_in_0_valid = io_in_2_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_RouteID = 16'h2; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_address = io_in_2_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_taskID = io_in_2_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 52:67]
  assign LockingRRArbiter_1_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_1_io_in_1_bits_address = 32'h0;
  assign LockingRRArbiter_1_io_in_1_bits_taskID = 10'h0;
  assign LockingRRArbiter_1_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_1_io_out_ready = LockingRRArbiter_2_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_clock = clock;
  assign LockingRRArbiter_2_io_in_0_valid = LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_0_bits_RouteID = LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_0_bits_address = LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_0_bits_taskID = LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_0_bits_Typ = LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_1_valid = LockingRRArbiter_1_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_1_bits_RouteID = LockingRRArbiter_1_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_1_bits_address = LockingRRArbiter_1_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_1_bits_taskID = LockingRRArbiter_1_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_in_1_bits_Typ = LockingRRArbiter_1_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_io_out_ready = io_out_ready; // @[ArbiterTree.scala 65:12]
endmodule
module RRArbiter_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  input  [31:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input  [31:0] io_in_1_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_data,
  output        io_chosen
);
  reg  _T_81; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  wire  _T_84; // @[Arbiter.scala 67:57]
  wire  _T_86; // @[Arbiter.scala 68:83]
  wire  _T_89; // @[Arbiter.scala 31:68]
  wire  _T_95; // @[Arbiter.scala 31:78]
  wire  _GEN_11; // @[Arbiter.scala 77:27]
  assign _T_84 = 1'h1 > _T_81; // @[Arbiter.scala 67:57]
  assign _T_86 = io_in_1_valid & _T_84; // @[Arbiter.scala 68:83]
  assign _T_89 = _T_86 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_95 = _T_89 == 1'h0; // @[Arbiter.scala 31:78]
  assign _GEN_11 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_86 == 1'h0; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_84 | _T_95; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_86 ? 1'h1 : _GEN_11; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_81 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_out_valid) begin
      _T_81 <= io_chosen;
    end
  end
endmodule
module Demux_3(
  input         io_en,
  input  [15:0] io_input_RouteID,
  input  [31:0] io_input_data,
  input         io_sel,
  output        io_outputs_0_valid,
  output [15:0] io_outputs_0_RouteID,
  output [31:0] io_outputs_0_data,
  output        io_outputs_1_valid,
  output [15:0] io_outputs_1_RouteID,
  output [31:0] io_outputs_1_data
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en ? _GEN_0 : 1'h0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_RouteID = io_input_RouteID; // @[Muxes.scala 23:19]
  assign io_outputs_0_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en ? io_sel : 1'h0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_RouteID = io_input_RouteID; // @[Muxes.scala 23:19]
  assign io_outputs_1_data = io_input_data; // @[Muxes.scala 23:19]
endmodule
module DeMuxTree_1(
  input         clock,
  input         reset,
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data,
  output        io_outputs_2_valid,
  output [31:0] io_outputs_2_data,
  input  [15:0] io_input_RouteID,
  input  [31:0] io_input_data,
  input         io_enable
);
  wire  Demux_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_1_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_1_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_1_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_1_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_1_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_1_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_1_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_2_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_2_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_2_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_2_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_2_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_2_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_2_io_outputs_1_data; // @[Muxes.scala 91:13]
  reg [15:0] _T_12_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_0;
  reg [31:0] _T_12_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_1;
  reg  _T_15; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_2;
  reg [15:0] _T_18_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_3;
  reg [31:0] _T_18_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_4;
  reg  _T_21; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_5;
  Demux_3 Demux ( // @[Muxes.scala 91:13]
    .io_en(Demux_io_en),
    .io_input_RouteID(Demux_io_input_RouteID),
    .io_input_data(Demux_io_input_data),
    .io_sel(Demux_io_sel),
    .io_outputs_0_valid(Demux_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_io_outputs_0_data),
    .io_outputs_1_valid(Demux_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_io_outputs_1_data)
  );
  Demux_3 Demux_1 ( // @[Muxes.scala 91:13]
    .io_en(Demux_1_io_en),
    .io_input_RouteID(Demux_1_io_input_RouteID),
    .io_input_data(Demux_1_io_input_data),
    .io_sel(Demux_1_io_sel),
    .io_outputs_0_valid(Demux_1_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_1_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_1_io_outputs_0_data),
    .io_outputs_1_valid(Demux_1_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_1_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_1_io_outputs_1_data)
  );
  Demux_3 Demux_2 ( // @[Muxes.scala 91:13]
    .io_en(Demux_2_io_en),
    .io_input_RouteID(Demux_2_io_input_RouteID),
    .io_input_data(Demux_2_io_input_data),
    .io_sel(Demux_2_io_sel),
    .io_outputs_0_valid(Demux_2_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_2_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_2_io_outputs_0_data),
    .io_outputs_1_valid(Demux_2_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_2_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_2_io_outputs_1_data)
  );
  assign io_outputs_0_valid = Demux_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_0_data = Demux_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_1_valid = Demux_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_1_data = Demux_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_2_valid = Demux_1_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_2_data = Demux_1_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign Demux_io_en = _T_15; // @[Muxes.scala 105:20]
  assign Demux_io_input_RouteID = _T_12_RouteID; // @[Muxes.scala 104:23]
  assign Demux_io_input_data = _T_12_data; // @[Muxes.scala 104:23]
  assign Demux_io_sel = _T_12_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_1_io_en = _T_21; // @[Muxes.scala 105:20]
  assign Demux_1_io_input_RouteID = _T_18_RouteID; // @[Muxes.scala 104:23]
  assign Demux_1_io_input_data = _T_18_data; // @[Muxes.scala 104:23]
  assign Demux_1_io_sel = _T_18_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_2_io_en = io_enable; // @[Muxes.scala 135:14]
  assign Demux_2_io_input_RouteID = io_input_RouteID; // @[Muxes.scala 134:17]
  assign Demux_2_io_input_data = io_input_data; // @[Muxes.scala 134:17]
  assign Demux_2_io_sel = io_input_RouteID[1]; // @[Muxes.scala 136:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12_RouteID = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_12_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_15 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_18_RouteID = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_18_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_21 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_12_RouteID <= Demux_2_io_outputs_0_RouteID;
    _T_12_data <= Demux_2_io_outputs_0_data;
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      _T_15 <= Demux_2_io_outputs_0_valid;
    end
    _T_18_RouteID <= Demux_2_io_outputs_1_RouteID;
    _T_18_data <= Demux_2_io_outputs_1_data;
    if (reset) begin
      _T_21 <= 1'h0;
    end else begin
      _T_21 <= Demux_2_io_outputs_1_valid;
    end
  end
endmodule
module ReadTableEntry(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [31:0] io_NodeReq_bits_address,
  input  [9:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_data,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output [31:0] io_output_bits_data,
  output        io_free
);
  reg  ID; // @[ReadMemoryController.scala 49:19]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_1;
  reg [31:0] request_R_address; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_2;
  reg [9:0] request_R_taskID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_3;
  reg [7:0] request_R_Typ; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_4;
  reg [63:0] bitmask; // @[ReadMemoryController.scala 56:29]
  reg [63:0] _RAND_5;
  reg [7:0] sendbytemask; // @[ReadMemoryController.scala 58:29]
  reg [31:0] _RAND_6;
  reg [31:0] ReqAddress; // @[ReadMemoryController.scala 62:27]
  reg [31:0] _RAND_7;
  reg  ptr; // @[ReadMemoryController.scala 66:27]
  reg [31:0] _RAND_8;
  reg [31:0] linebuffer_0; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_9;
  reg [31:0] linebuffer_1; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[ReadMemoryController.scala 73:68]
  reg [31:0] _RAND_11;
  wire [2:0] _T_100; // @[Cat.scala 30:58]
  wire [31:0] _GEN_57; // @[ReadMemoryController.scala 96:37]
  wire [32:0] _T_101; // @[ReadMemoryController.scala 96:37]
  reg  isWrite; // @[ReadMemoryController.scala 100:24]
  reg [31:0] _RAND_12;
  wire  _T_109; // @[Decoupled.scala 37:37]
  wire [29:0] _T_110; // @[ReadMemoryController.scala 115:44]
  wire [31:0] _GEN_58; // @[ReadMemoryController.scala 115:69]
  wire [31:0] _T_111; // @[ReadMemoryController.scala 115:69]
  wire  _T_112; // @[helpers.scala 27:24]
  wire  _T_113; // @[helpers.scala 27:47]
  wire  _T_114; // @[helpers.scala 27:40]
  wire  _T_120; // @[helpers.scala 28:15]
  wire  _T_121; // @[helpers.scala 28:38]
  wire  _T_122; // @[helpers.scala 28:31]
  wire  _T_128; // @[helpers.scala 29:17]
  wire  _T_129; // @[helpers.scala 29:40]
  wire  _T_130; // @[helpers.scala 29:33]
  wire [63:0] _T_141; // @[helpers.scala 29:12]
  wire [63:0] _T_142; // @[helpers.scala 28:10]
  wire [63:0] _T_143; // @[helpers.scala 27:19]
  wire [1:0] _T_144; // @[helpers.scala 39:32]
  wire [4:0] _T_146; // @[Cat.scala 30:58]
  wire [94:0] _GEN_59; // @[helpers.scala 40:26]
  wire [94:0] _T_147; // @[helpers.scala 40:26]
  wire [7:0] _T_173; // @[helpers.scala 50:12]
  wire [7:0] _T_174; // @[helpers.scala 49:10]
  wire [7:0] _T_175; // @[helpers.scala 48:19]
  wire [10:0] _GEN_60; // @[helpers.scala 20:26]
  wire [10:0] _T_177; // @[helpers.scala 20:26]
  wire [7:0] _GEN_0; // @[ReadMemoryController.scala 111:28]
  wire [9:0] _GEN_1; // @[ReadMemoryController.scala 111:28]
  wire [31:0] _GEN_2; // @[ReadMemoryController.scala 111:28]
  wire [15:0] _GEN_3; // @[ReadMemoryController.scala 111:28]
  wire [31:0] _GEN_4; // @[ReadMemoryController.scala 111:28]
  wire [94:0] _GEN_5; // @[ReadMemoryController.scala 111:28]
  wire [10:0] _GEN_6; // @[ReadMemoryController.scala 111:28]
  wire  _T_178; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_7; // @[ReadMemoryController.scala 135:32]
  wire  _T_180; // @[Conditional.scala 37:30]
  wire [3:0] _T_182; // @[ReadMemoryController.scala 144:38]
  wire [10:0] _GEN_8; // @[ReadMemoryController.scala 142:29]
  wire [1:0] _GEN_9; // @[ReadMemoryController.scala 142:29]
  wire  _T_183; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_10; // @[ReadMemoryController.scala 152:25]
  wire [31:0] _GEN_11; // @[ReadMemoryController.scala 152:25]
  wire [1:0] _T_188; // @[ReadMemoryController.scala 154:20]
  wire  _T_189; // @[ReadMemoryController.scala 154:20]
  wire  _T_191; // @[ReadMemoryController.scala 156:27]
  wire [1:0] _GEN_12; // @[ReadMemoryController.scala 156:55]
  wire [31:0] _GEN_13; // @[ReadMemoryController.scala 150:30]
  wire [31:0] _GEN_14; // @[ReadMemoryController.scala 150:30]
  wire  _GEN_15; // @[ReadMemoryController.scala 150:30]
  wire [1:0] _GEN_16; // @[ReadMemoryController.scala 150:30]
  wire  _T_192; // @[Conditional.scala 37:30]
  wire [63:0] _T_194; // @[ReadMemoryController.scala 165:29]
  wire [63:0] _T_195; // @[ReadMemoryController.scala 165:36]
  wire [1:0] _T_196; // @[ReadMemoryController.scala 165:71]
  wire [4:0] _T_198; // @[Cat.scala 30:58]
  wire [63:0] _T_199; // @[ReadMemoryController.scala 165:47]
  wire  _T_200; // @[helpers.scala 63:30]
  wire [63:0] _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_53; // @[Conditional.scala 40:58]
  wire [31:0] output$; // @[ReadMemoryController.scala 165:14]
  wire  _T_201; // @[helpers.scala 63:57]
  wire [15:0] _T_205; // @[Bitwise.scala 72:12]
  wire [15:0] _T_206; // @[helpers.scala 63:68]
  wire [31:0] _T_207; // @[Cat.scala 30:58]
  wire  _T_208; // @[helpers.scala 64:22]
  wire [31:0] _T_215; // @[Cat.scala 30:58]
  wire  _T_216; // @[helpers.scala 65:24]
  wire  _T_217; // @[helpers.scala 65:51]
  wire [23:0] _T_221; // @[Bitwise.scala 72:12]
  wire [7:0] _T_222; // @[helpers.scala 65:61]
  wire [31:0] _T_223; // @[Cat.scala 30:58]
  wire  _T_224; // @[helpers.scala 66:26]
  wire [31:0] _T_231; // @[Cat.scala 30:58]
  wire [31:0] _T_233; // @[helpers.scala 66:14]
  wire [31:0] _T_234; // @[helpers.scala 65:12]
  wire [31:0] _T_235; // @[helpers.scala 64:10]
  wire [31:0] _T_236; // @[helpers.scala 63:18]
  wire [1:0] _GEN_17; // @[ReadMemoryController.scala 176:29]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_23; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_24; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_27; // @[Conditional.scala 39:67]
  wire  _GEN_28; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_36; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_37; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_38; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_46; // @[Conditional.scala 40:58]
  wire [10:0] _GEN_48; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_49; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  assign _T_100 = {ptr,2'h0}; // @[Cat.scala 30:58]
  assign _GEN_57 = {{29'd0}, _T_100}; // @[ReadMemoryController.scala 96:37]
  assign _T_101 = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:37]
  assign _T_109 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 37:37]
  assign _T_110 = io_NodeReq_bits_address[31:2]; // @[ReadMemoryController.scala 115:44]
  assign _GEN_58 = {{2'd0}, _T_110}; // @[ReadMemoryController.scala 115:69]
  assign _T_111 = _GEN_58 << 2; // @[ReadMemoryController.scala 115:69]
  assign _T_112 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_113 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_114 = _T_112 | _T_113; // @[helpers.scala 27:40]
  assign _T_120 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_121 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_122 = _T_120 | _T_121; // @[helpers.scala 28:31]
  assign _T_128 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_129 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_130 = _T_128 | _T_129; // @[helpers.scala 29:33]
  assign _T_141 = _T_130 ? 64'hffffffff : 64'hffffffffffffffff; // @[helpers.scala 29:12]
  assign _T_142 = _T_122 ? 64'hff : _T_141; // @[helpers.scala 28:10]
  assign _T_143 = _T_114 ? 64'hffff : _T_142; // @[helpers.scala 27:19]
  assign _T_144 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_146 = {_T_144,3'h0}; // @[Cat.scala 30:58]
  assign _GEN_59 = {{31'd0}, _T_143}; // @[helpers.scala 40:26]
  assign _T_147 = _GEN_59 << _T_146; // @[helpers.scala 40:26]
  assign _T_173 = _T_130 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_174 = _T_122 ? 8'h1 : _T_173; // @[helpers.scala 49:10]
  assign _T_175 = _T_114 ? 8'h3 : _T_174; // @[helpers.scala 48:19]
  assign _GEN_60 = {{3'd0}, _T_175}; // @[helpers.scala 20:26]
  assign _T_177 = _GEN_60 << _T_144; // @[helpers.scala 20:26]
  assign _GEN_0 = _T_109 ? io_NodeReq_bits_Typ : request_R_Typ; // @[ReadMemoryController.scala 111:28]
  assign _GEN_1 = _T_109 ? io_NodeReq_bits_taskID : request_R_taskID; // @[ReadMemoryController.scala 111:28]
  assign _GEN_2 = _T_109 ? io_NodeReq_bits_address : request_R_address; // @[ReadMemoryController.scala 111:28]
  assign _GEN_3 = _T_109 ? io_NodeReq_bits_RouteID : request_R_RouteID; // @[ReadMemoryController.scala 111:28]
  assign _GEN_4 = _T_109 ? _T_111 : ReqAddress; // @[ReadMemoryController.scala 111:28]
  assign _GEN_5 = _T_109 ? _T_147 : {{31'd0}, bitmask}; // @[ReadMemoryController.scala 111:28]
  assign _GEN_6 = _T_109 ? _T_177 : {{3'd0}, sendbytemask}; // @[ReadMemoryController.scala 111:28]
  assign _T_178 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_7 = _T_109 ? 2'h1 : state; // @[ReadMemoryController.scala 135:32]
  assign _T_180 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_182 = sendbytemask[7:4]; // @[ReadMemoryController.scala 144:38]
  assign _GEN_8 = io_MemReq_ready ? {{7'd0}, _T_182} : _GEN_6; // @[ReadMemoryController.scala 142:29]
  assign _GEN_9 = io_MemReq_ready ? 2'h2 : state; // @[ReadMemoryController.scala 142:29]
  assign _T_183 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_10 = 1'h0 == ptr ? io_MemResp_data : linebuffer_0; // @[ReadMemoryController.scala 152:25]
  assign _GEN_11 = ptr ? io_MemResp_data : linebuffer_1; // @[ReadMemoryController.scala 152:25]
  assign _T_188 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_189 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_191 = sendbytemask == 8'h0; // @[ReadMemoryController.scala 156:27]
  assign _GEN_12 = _T_191 ? 2'h3 : 2'h1; // @[ReadMemoryController.scala 156:55]
  assign _GEN_13 = io_MemResp_valid ? _GEN_10 : linebuffer_0; // @[ReadMemoryController.scala 150:30]
  assign _GEN_14 = io_MemResp_valid ? _GEN_11 : linebuffer_1; // @[ReadMemoryController.scala 150:30]
  assign _GEN_15 = io_MemResp_valid ? _T_189 : ptr; // @[ReadMemoryController.scala 150:30]
  assign _GEN_16 = io_MemResp_valid ? _GEN_12 : state; // @[ReadMemoryController.scala 150:30]
  assign _T_192 = 2'h3 == state; // @[Conditional.scala 37:30]
  assign _T_194 = {linebuffer_1,linebuffer_0}; // @[ReadMemoryController.scala 165:29]
  assign _T_195 = _T_194 & bitmask; // @[ReadMemoryController.scala 165:36]
  assign _T_196 = request_R_address[1:0]; // @[ReadMemoryController.scala 165:71]
  assign _T_198 = {_T_196,3'h0}; // @[Cat.scala 30:58]
  assign _T_199 = _T_195 >> _T_198; // @[ReadMemoryController.scala 165:47]
  assign _T_200 = request_R_Typ == 8'h2; // @[helpers.scala 63:30]
  assign _GEN_20 = _T_192 ? _T_199 : 64'h0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_183 ? 64'h0 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_180 ? 64'h0 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_178 ? 64'h0 : _GEN_42; // @[Conditional.scala 40:58]
  assign output$ = _GEN_53[31:0]; // @[ReadMemoryController.scala 165:14]
  assign _T_201 = output$[15]; // @[helpers.scala 63:57]
  assign _T_205 = _T_201 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  assign _T_206 = output$[15:0]; // @[helpers.scala 63:68]
  assign _T_207 = {_T_205,_T_206}; // @[Cat.scala 30:58]
  assign _T_208 = request_R_Typ == 8'h6; // @[helpers.scala 64:22]
  assign _T_215 = {16'h0,_T_206}; // @[Cat.scala 30:58]
  assign _T_216 = request_R_Typ == 8'h1; // @[helpers.scala 65:24]
  assign _T_217 = output$[7]; // @[helpers.scala 65:51]
  assign _T_221 = _T_217 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_222 = output$[7:0]; // @[helpers.scala 65:61]
  assign _T_223 = {_T_221,_T_222}; // @[Cat.scala 30:58]
  assign _T_224 = request_R_Typ == 8'h5; // @[helpers.scala 66:26]
  assign _T_231 = {24'h0,_T_222}; // @[Cat.scala 30:58]
  assign _T_233 = _T_224 ? _T_231 : output$; // @[helpers.scala 66:14]
  assign _T_234 = _T_216 ? _T_223 : _T_233; // @[helpers.scala 65:12]
  assign _T_235 = _T_208 ? _T_215 : _T_234; // @[helpers.scala 64:10]
  assign _T_236 = _T_200 ? _T_207 : _T_235; // @[helpers.scala 63:18]
  assign _GEN_17 = io_output_ready ? 2'h0 : state; // @[ReadMemoryController.scala 176:29]
  assign _GEN_21 = _T_192 ? _T_236 : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_23 = _T_192 ? 1'h0 : ptr; // @[Conditional.scala 39:67]
  assign _GEN_24 = _T_192 ? _GEN_17 : state; // @[Conditional.scala 39:67]
  assign _GEN_26 = _T_183 ? _GEN_13 : linebuffer_0; // @[Conditional.scala 39:67]
  assign _GEN_27 = _T_183 ? _GEN_14 : linebuffer_1; // @[Conditional.scala 39:67]
  assign _GEN_28 = _T_183 ? _GEN_15 : _GEN_23; // @[Conditional.scala 39:67]
  assign _GEN_29 = _T_183 ? _GEN_16 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_183 ? 1'h0 : _T_192; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_183 ? 32'h0 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_180 ? _GEN_8 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_180 ? _GEN_9 : _GEN_29; // @[Conditional.scala 39:67]
  assign _GEN_38 = _T_180 ? linebuffer_0 : _GEN_26; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_180 ? linebuffer_1 : _GEN_27; // @[Conditional.scala 39:67]
  assign _GEN_40 = _T_180 ? ptr : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_180 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_180 ? 32'h0 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_46 = _T_178 ? _GEN_7 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_178 ? _GEN_6 : _GEN_36; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_178 ? linebuffer_0 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_178 ? linebuffer_1 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_178 ? ptr : _GEN_40; // @[Conditional.scala 40:58]
  assign io_NodeReq_ready = state == 2'h0; // @[ReadMemoryController.scala 83:20]
  assign io_MemReq_valid = _T_178 ? 1'h0 : _T_180; // @[ReadMemoryController.scala 95:19 ReadMemoryController.scala 140:23]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:23]
  assign io_MemReq_bits_tag = {{7'd0}, ID}; // @[ReadMemoryController.scala 99:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[ReadMemoryController.scala 104:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[ReadMemoryController.scala 101:26]
  assign io_output_valid = _T_178 ? 1'h0 : _GEN_41; // @[ReadMemoryController.scala 90:19 ReadMemoryController.scala 164:23]
  assign io_output_bits_RouteID = request_R_RouteID; // @[ReadMemoryController.scala 91:26]
  assign io_output_bits_data = _T_178 ? 32'h0 : _GEN_43; // @[ReadMemoryController.scala 93:23 ReadMemoryController.scala 168:29]
  assign io_free = state == 2'h0; // @[ReadMemoryController.scala 81:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_address = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_R_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  request_R_Typ = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  bitmask = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sendbytemask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ReqAddress = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ptr = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  linebuffer_0 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  linebuffer_1 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  isWrite = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    ID <= reset;
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_109) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_address <= 32'h0;
    end else begin
      if (_T_109) begin
        request_R_address <= io_NodeReq_bits_address;
      end
    end
    if (reset) begin
      request_R_taskID <= 10'h0;
    end else begin
      if (_T_109) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      request_R_Typ <= 8'h3;
    end else begin
      if (_T_109) begin
        request_R_Typ <= io_NodeReq_bits_Typ;
      end
    end
    if (reset) begin
      bitmask <= 64'h0;
    end else begin
      bitmask <= _GEN_5[63:0];
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_48[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_109) begin
        ReqAddress <= _T_111;
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (!(_T_178)) begin
        if (!(_T_180)) begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              ptr <= _T_189;
            end
          end else begin
            if (_T_192) begin
              ptr <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (!(_T_178)) begin
        if (!(_T_180)) begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              if (1'h0 == ptr) begin
                linebuffer_0 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (!(_T_178)) begin
        if (!(_T_180)) begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              if (ptr) begin
                linebuffer_1 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_178) begin
        if (_T_109) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_180) begin
          if (io_MemReq_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              if (_T_191) begin
                state <= 2'h3;
              end else begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_192) begin
              if (io_output_ready) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    isWrite <= reset;
  end
endmodule
module ReadTableEntry_1(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [31:0] io_NodeReq_bits_address,
  input  [9:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_data,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output [31:0] io_output_bits_data,
  output        io_free
);
  reg  ID; // @[ReadMemoryController.scala 49:19]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_1;
  reg [31:0] request_R_address; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_2;
  reg [9:0] request_R_taskID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_3;
  reg [7:0] request_R_Typ; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_4;
  reg [63:0] bitmask; // @[ReadMemoryController.scala 56:29]
  reg [63:0] _RAND_5;
  reg [7:0] sendbytemask; // @[ReadMemoryController.scala 58:29]
  reg [31:0] _RAND_6;
  reg [31:0] ReqAddress; // @[ReadMemoryController.scala 62:27]
  reg [31:0] _RAND_7;
  reg  ptr; // @[ReadMemoryController.scala 66:27]
  reg [31:0] _RAND_8;
  reg [31:0] linebuffer_0; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_9;
  reg [31:0] linebuffer_1; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[ReadMemoryController.scala 73:68]
  reg [31:0] _RAND_11;
  wire [2:0] _T_100; // @[Cat.scala 30:58]
  wire [31:0] _GEN_57; // @[ReadMemoryController.scala 96:37]
  wire [32:0] _T_101; // @[ReadMemoryController.scala 96:37]
  reg  isWrite; // @[ReadMemoryController.scala 100:24]
  reg [31:0] _RAND_12;
  wire  _T_109; // @[Decoupled.scala 37:37]
  wire [29:0] _T_110; // @[ReadMemoryController.scala 115:44]
  wire [31:0] _GEN_58; // @[ReadMemoryController.scala 115:69]
  wire [31:0] _T_111; // @[ReadMemoryController.scala 115:69]
  wire  _T_112; // @[helpers.scala 27:24]
  wire  _T_113; // @[helpers.scala 27:47]
  wire  _T_114; // @[helpers.scala 27:40]
  wire  _T_120; // @[helpers.scala 28:15]
  wire  _T_121; // @[helpers.scala 28:38]
  wire  _T_122; // @[helpers.scala 28:31]
  wire  _T_128; // @[helpers.scala 29:17]
  wire  _T_129; // @[helpers.scala 29:40]
  wire  _T_130; // @[helpers.scala 29:33]
  wire [63:0] _T_141; // @[helpers.scala 29:12]
  wire [63:0] _T_142; // @[helpers.scala 28:10]
  wire [63:0] _T_143; // @[helpers.scala 27:19]
  wire [1:0] _T_144; // @[helpers.scala 39:32]
  wire [4:0] _T_146; // @[Cat.scala 30:58]
  wire [94:0] _GEN_59; // @[helpers.scala 40:26]
  wire [94:0] _T_147; // @[helpers.scala 40:26]
  wire [7:0] _T_173; // @[helpers.scala 50:12]
  wire [7:0] _T_174; // @[helpers.scala 49:10]
  wire [7:0] _T_175; // @[helpers.scala 48:19]
  wire [10:0] _GEN_60; // @[helpers.scala 20:26]
  wire [10:0] _T_177; // @[helpers.scala 20:26]
  wire [7:0] _GEN_0; // @[ReadMemoryController.scala 111:28]
  wire [9:0] _GEN_1; // @[ReadMemoryController.scala 111:28]
  wire [31:0] _GEN_2; // @[ReadMemoryController.scala 111:28]
  wire [15:0] _GEN_3; // @[ReadMemoryController.scala 111:28]
  wire [31:0] _GEN_4; // @[ReadMemoryController.scala 111:28]
  wire [94:0] _GEN_5; // @[ReadMemoryController.scala 111:28]
  wire [10:0] _GEN_6; // @[ReadMemoryController.scala 111:28]
  wire  _T_178; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_7; // @[ReadMemoryController.scala 135:32]
  wire  _T_180; // @[Conditional.scala 37:30]
  wire [3:0] _T_182; // @[ReadMemoryController.scala 144:38]
  wire [10:0] _GEN_8; // @[ReadMemoryController.scala 142:29]
  wire [1:0] _GEN_9; // @[ReadMemoryController.scala 142:29]
  wire  _T_183; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_10; // @[ReadMemoryController.scala 152:25]
  wire [31:0] _GEN_11; // @[ReadMemoryController.scala 152:25]
  wire [1:0] _T_188; // @[ReadMemoryController.scala 154:20]
  wire  _T_189; // @[ReadMemoryController.scala 154:20]
  wire  _T_191; // @[ReadMemoryController.scala 156:27]
  wire [1:0] _GEN_12; // @[ReadMemoryController.scala 156:55]
  wire [31:0] _GEN_13; // @[ReadMemoryController.scala 150:30]
  wire [31:0] _GEN_14; // @[ReadMemoryController.scala 150:30]
  wire  _GEN_15; // @[ReadMemoryController.scala 150:30]
  wire [1:0] _GEN_16; // @[ReadMemoryController.scala 150:30]
  wire  _T_192; // @[Conditional.scala 37:30]
  wire [63:0] _T_194; // @[ReadMemoryController.scala 165:29]
  wire [63:0] _T_195; // @[ReadMemoryController.scala 165:36]
  wire [1:0] _T_196; // @[ReadMemoryController.scala 165:71]
  wire [4:0] _T_198; // @[Cat.scala 30:58]
  wire [63:0] _T_199; // @[ReadMemoryController.scala 165:47]
  wire  _T_200; // @[helpers.scala 63:30]
  wire [63:0] _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_53; // @[Conditional.scala 40:58]
  wire [31:0] output$; // @[ReadMemoryController.scala 165:14]
  wire  _T_201; // @[helpers.scala 63:57]
  wire [15:0] _T_205; // @[Bitwise.scala 72:12]
  wire [15:0] _T_206; // @[helpers.scala 63:68]
  wire [31:0] _T_207; // @[Cat.scala 30:58]
  wire  _T_208; // @[helpers.scala 64:22]
  wire [31:0] _T_215; // @[Cat.scala 30:58]
  wire  _T_216; // @[helpers.scala 65:24]
  wire  _T_217; // @[helpers.scala 65:51]
  wire [23:0] _T_221; // @[Bitwise.scala 72:12]
  wire [7:0] _T_222; // @[helpers.scala 65:61]
  wire [31:0] _T_223; // @[Cat.scala 30:58]
  wire  _T_224; // @[helpers.scala 66:26]
  wire [31:0] _T_231; // @[Cat.scala 30:58]
  wire [31:0] _T_233; // @[helpers.scala 66:14]
  wire [31:0] _T_234; // @[helpers.scala 65:12]
  wire [31:0] _T_235; // @[helpers.scala 64:10]
  wire [31:0] _T_236; // @[helpers.scala 63:18]
  wire [1:0] _GEN_17; // @[ReadMemoryController.scala 176:29]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_23; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_24; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_26; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_27; // @[Conditional.scala 39:67]
  wire  _GEN_28; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_36; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_37; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_38; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_46; // @[Conditional.scala 40:58]
  wire [10:0] _GEN_48; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_49; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  assign _T_100 = {ptr,2'h0}; // @[Cat.scala 30:58]
  assign _GEN_57 = {{29'd0}, _T_100}; // @[ReadMemoryController.scala 96:37]
  assign _T_101 = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:37]
  assign _T_109 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 37:37]
  assign _T_110 = io_NodeReq_bits_address[31:2]; // @[ReadMemoryController.scala 115:44]
  assign _GEN_58 = {{2'd0}, _T_110}; // @[ReadMemoryController.scala 115:69]
  assign _T_111 = _GEN_58 << 2; // @[ReadMemoryController.scala 115:69]
  assign _T_112 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_113 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_114 = _T_112 | _T_113; // @[helpers.scala 27:40]
  assign _T_120 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_121 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_122 = _T_120 | _T_121; // @[helpers.scala 28:31]
  assign _T_128 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_129 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_130 = _T_128 | _T_129; // @[helpers.scala 29:33]
  assign _T_141 = _T_130 ? 64'hffffffff : 64'hffffffffffffffff; // @[helpers.scala 29:12]
  assign _T_142 = _T_122 ? 64'hff : _T_141; // @[helpers.scala 28:10]
  assign _T_143 = _T_114 ? 64'hffff : _T_142; // @[helpers.scala 27:19]
  assign _T_144 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_146 = {_T_144,3'h0}; // @[Cat.scala 30:58]
  assign _GEN_59 = {{31'd0}, _T_143}; // @[helpers.scala 40:26]
  assign _T_147 = _GEN_59 << _T_146; // @[helpers.scala 40:26]
  assign _T_173 = _T_130 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_174 = _T_122 ? 8'h1 : _T_173; // @[helpers.scala 49:10]
  assign _T_175 = _T_114 ? 8'h3 : _T_174; // @[helpers.scala 48:19]
  assign _GEN_60 = {{3'd0}, _T_175}; // @[helpers.scala 20:26]
  assign _T_177 = _GEN_60 << _T_144; // @[helpers.scala 20:26]
  assign _GEN_0 = _T_109 ? io_NodeReq_bits_Typ : request_R_Typ; // @[ReadMemoryController.scala 111:28]
  assign _GEN_1 = _T_109 ? io_NodeReq_bits_taskID : request_R_taskID; // @[ReadMemoryController.scala 111:28]
  assign _GEN_2 = _T_109 ? io_NodeReq_bits_address : request_R_address; // @[ReadMemoryController.scala 111:28]
  assign _GEN_3 = _T_109 ? io_NodeReq_bits_RouteID : request_R_RouteID; // @[ReadMemoryController.scala 111:28]
  assign _GEN_4 = _T_109 ? _T_111 : ReqAddress; // @[ReadMemoryController.scala 111:28]
  assign _GEN_5 = _T_109 ? _T_147 : {{31'd0}, bitmask}; // @[ReadMemoryController.scala 111:28]
  assign _GEN_6 = _T_109 ? _T_177 : {{3'd0}, sendbytemask}; // @[ReadMemoryController.scala 111:28]
  assign _T_178 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_7 = _T_109 ? 2'h1 : state; // @[ReadMemoryController.scala 135:32]
  assign _T_180 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_182 = sendbytemask[7:4]; // @[ReadMemoryController.scala 144:38]
  assign _GEN_8 = io_MemReq_ready ? {{7'd0}, _T_182} : _GEN_6; // @[ReadMemoryController.scala 142:29]
  assign _GEN_9 = io_MemReq_ready ? 2'h2 : state; // @[ReadMemoryController.scala 142:29]
  assign _T_183 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_10 = 1'h0 == ptr ? io_MemResp_data : linebuffer_0; // @[ReadMemoryController.scala 152:25]
  assign _GEN_11 = ptr ? io_MemResp_data : linebuffer_1; // @[ReadMemoryController.scala 152:25]
  assign _T_188 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_189 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_191 = sendbytemask == 8'h0; // @[ReadMemoryController.scala 156:27]
  assign _GEN_12 = _T_191 ? 2'h3 : 2'h1; // @[ReadMemoryController.scala 156:55]
  assign _GEN_13 = io_MemResp_valid ? _GEN_10 : linebuffer_0; // @[ReadMemoryController.scala 150:30]
  assign _GEN_14 = io_MemResp_valid ? _GEN_11 : linebuffer_1; // @[ReadMemoryController.scala 150:30]
  assign _GEN_15 = io_MemResp_valid ? _T_189 : ptr; // @[ReadMemoryController.scala 150:30]
  assign _GEN_16 = io_MemResp_valid ? _GEN_12 : state; // @[ReadMemoryController.scala 150:30]
  assign _T_192 = 2'h3 == state; // @[Conditional.scala 37:30]
  assign _T_194 = {linebuffer_1,linebuffer_0}; // @[ReadMemoryController.scala 165:29]
  assign _T_195 = _T_194 & bitmask; // @[ReadMemoryController.scala 165:36]
  assign _T_196 = request_R_address[1:0]; // @[ReadMemoryController.scala 165:71]
  assign _T_198 = {_T_196,3'h0}; // @[Cat.scala 30:58]
  assign _T_199 = _T_195 >> _T_198; // @[ReadMemoryController.scala 165:47]
  assign _T_200 = request_R_Typ == 8'h2; // @[helpers.scala 63:30]
  assign _GEN_20 = _T_192 ? _T_199 : 64'h0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_183 ? 64'h0 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_180 ? 64'h0 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_178 ? 64'h0 : _GEN_42; // @[Conditional.scala 40:58]
  assign output$ = _GEN_53[31:0]; // @[ReadMemoryController.scala 165:14]
  assign _T_201 = output$[15]; // @[helpers.scala 63:57]
  assign _T_205 = _T_201 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  assign _T_206 = output$[15:0]; // @[helpers.scala 63:68]
  assign _T_207 = {_T_205,_T_206}; // @[Cat.scala 30:58]
  assign _T_208 = request_R_Typ == 8'h6; // @[helpers.scala 64:22]
  assign _T_215 = {16'h0,_T_206}; // @[Cat.scala 30:58]
  assign _T_216 = request_R_Typ == 8'h1; // @[helpers.scala 65:24]
  assign _T_217 = output$[7]; // @[helpers.scala 65:51]
  assign _T_221 = _T_217 ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  assign _T_222 = output$[7:0]; // @[helpers.scala 65:61]
  assign _T_223 = {_T_221,_T_222}; // @[Cat.scala 30:58]
  assign _T_224 = request_R_Typ == 8'h5; // @[helpers.scala 66:26]
  assign _T_231 = {24'h0,_T_222}; // @[Cat.scala 30:58]
  assign _T_233 = _T_224 ? _T_231 : output$; // @[helpers.scala 66:14]
  assign _T_234 = _T_216 ? _T_223 : _T_233; // @[helpers.scala 65:12]
  assign _T_235 = _T_208 ? _T_215 : _T_234; // @[helpers.scala 64:10]
  assign _T_236 = _T_200 ? _T_207 : _T_235; // @[helpers.scala 63:18]
  assign _GEN_17 = io_output_ready ? 2'h0 : state; // @[ReadMemoryController.scala 176:29]
  assign _GEN_21 = _T_192 ? _T_236 : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_23 = _T_192 ? 1'h0 : ptr; // @[Conditional.scala 39:67]
  assign _GEN_24 = _T_192 ? _GEN_17 : state; // @[Conditional.scala 39:67]
  assign _GEN_26 = _T_183 ? _GEN_13 : linebuffer_0; // @[Conditional.scala 39:67]
  assign _GEN_27 = _T_183 ? _GEN_14 : linebuffer_1; // @[Conditional.scala 39:67]
  assign _GEN_28 = _T_183 ? _GEN_15 : _GEN_23; // @[Conditional.scala 39:67]
  assign _GEN_29 = _T_183 ? _GEN_16 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_183 ? 1'h0 : _T_192; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_183 ? 32'h0 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_180 ? _GEN_8 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_180 ? _GEN_9 : _GEN_29; // @[Conditional.scala 39:67]
  assign _GEN_38 = _T_180 ? linebuffer_0 : _GEN_26; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_180 ? linebuffer_1 : _GEN_27; // @[Conditional.scala 39:67]
  assign _GEN_40 = _T_180 ? ptr : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_180 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_180 ? 32'h0 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_46 = _T_178 ? _GEN_7 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_178 ? _GEN_6 : _GEN_36; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_178 ? linebuffer_0 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_178 ? linebuffer_1 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_178 ? ptr : _GEN_40; // @[Conditional.scala 40:58]
  assign io_NodeReq_ready = state == 2'h0; // @[ReadMemoryController.scala 83:20]
  assign io_MemReq_valid = _T_178 ? 1'h0 : _T_180; // @[ReadMemoryController.scala 95:19 ReadMemoryController.scala 140:23]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:23]
  assign io_MemReq_bits_tag = {{7'd0}, ID}; // @[ReadMemoryController.scala 99:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[ReadMemoryController.scala 104:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[ReadMemoryController.scala 101:26]
  assign io_output_valid = _T_178 ? 1'h0 : _GEN_41; // @[ReadMemoryController.scala 90:19 ReadMemoryController.scala 164:23]
  assign io_output_bits_RouteID = request_R_RouteID; // @[ReadMemoryController.scala 91:26]
  assign io_output_bits_data = _T_178 ? 32'h0 : _GEN_43; // @[ReadMemoryController.scala 93:23 ReadMemoryController.scala 168:29]
  assign io_free = state == 2'h0; // @[ReadMemoryController.scala 81:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_address = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_R_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  request_R_Typ = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  bitmask = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sendbytemask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ReqAddress = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ptr = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  linebuffer_0 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  linebuffer_1 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  isWrite = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ID <= 1'h0;
    end else begin
      ID <= 1'h1;
    end
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_109) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_address <= 32'h0;
    end else begin
      if (_T_109) begin
        request_R_address <= io_NodeReq_bits_address;
      end
    end
    if (reset) begin
      request_R_taskID <= 10'h0;
    end else begin
      if (_T_109) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      request_R_Typ <= 8'h3;
    end else begin
      if (_T_109) begin
        request_R_Typ <= io_NodeReq_bits_Typ;
      end
    end
    if (reset) begin
      bitmask <= 64'h0;
    end else begin
      bitmask <= _GEN_5[63:0];
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_48[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_109) begin
        ReqAddress <= _T_111;
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (!(_T_178)) begin
        if (!(_T_180)) begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              ptr <= _T_189;
            end
          end else begin
            if (_T_192) begin
              ptr <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (!(_T_178)) begin
        if (!(_T_180)) begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              if (1'h0 == ptr) begin
                linebuffer_0 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (!(_T_178)) begin
        if (!(_T_180)) begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              if (ptr) begin
                linebuffer_1 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_178) begin
        if (_T_109) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_180) begin
          if (io_MemReq_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_183) begin
            if (io_MemResp_valid) begin
              if (_T_191) begin
                state <= 2'h3;
              end else begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_192) begin
              if (io_output_ready) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    isWrite <= reset;
  end
endmodule
module ReadMemoryController(
  input         clock,
  input         reset,
  output        io_ReadIn_0_ready,
  input         io_ReadIn_0_valid,
  input  [31:0] io_ReadIn_0_bits_address,
  input  [9:0]  io_ReadIn_0_bits_taskID,
  output        io_ReadIn_1_ready,
  input         io_ReadIn_1_valid,
  input  [31:0] io_ReadIn_1_bits_address,
  input  [9:0]  io_ReadIn_1_bits_taskID,
  output        io_ReadIn_2_ready,
  input         io_ReadIn_2_valid,
  input  [31:0] io_ReadIn_2_bits_address,
  input  [9:0]  io_ReadIn_2_bits_taskID,
  output        io_ReadOut_0_valid,
  output [31:0] io_ReadOut_0_data,
  output        io_ReadOut_1_valid,
  output [31:0] io_ReadOut_1_data,
  output        io_ReadOut_2_valid,
  output [31:0] io_ReadOut_2_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag
);
  wire  in_arb_clock; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_0_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_0_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_0_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [9:0] in_arb_io_in_0_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_1_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_1_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_1_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [9:0] in_arb_io_in_1_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_2_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_2_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_2_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [9:0] in_arb_io_in_2_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_out_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_out_valid; // @[ReadMemoryController.scala 221:25]
  wire [15:0] in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_out_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [9:0] in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire [7:0] in_arb_io_out_bits_Typ; // @[ReadMemoryController.scala 221:25]
  wire  alloc_arb_io_in_0_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_0_valid; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_1_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_1_valid; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_out_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_out_valid; // @[ReadMemoryController.scala 223:25]
  wire  cachereq_arb_io_in_0_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_0_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [9:0] cachereq_arb_io_in_0_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [9:0] cachereq_arb_io_in_1_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [9:0] cachereq_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cacheresp_demux_io_en; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_sel; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[ReadMemoryController.scala 228:31]
  wire  out_arb_clock; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_0_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_0_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_in_0_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_in_0_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_1_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_1_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_in_1_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_in_1_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_out_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_out_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_out_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_chosen; // @[ReadMemoryController.scala 231:25]
  wire  out_demux_clock; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_reset; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_0_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_1_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_2_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_2_data; // @[ReadMemoryController.scala 232:25]
  wire [15:0] out_demux_io_input_RouteID; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_input_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_enable; // @[ReadMemoryController.scala 232:25]
  wire  ReadTable_0_clock; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_reset; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_NodeReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_NodeReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_0_io_NodeReq_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_NodeReq_bits_address; // @[ReadMemoryController.scala 251:28]
  wire [9:0] ReadTable_0_io_NodeReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_0_io_NodeReq_bits_Typ; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_MemReq_bits_addr; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_0_io_MemReq_bits_tag; // @[ReadMemoryController.scala 251:28]
  wire [9:0] ReadTable_0_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemResp_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_MemResp_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_output_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_output_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_0_io_output_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_output_bits_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_free; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_clock; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_reset; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_NodeReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_NodeReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_1_io_NodeReq_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_NodeReq_bits_address; // @[ReadMemoryController.scala 251:28]
  wire [9:0] ReadTable_1_io_NodeReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_1_io_NodeReq_bits_Typ; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_MemReq_bits_addr; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_1_io_MemReq_bits_tag; // @[ReadMemoryController.scala 251:28]
  wire [9:0] ReadTable_1_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemResp_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_MemResp_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_output_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_output_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_1_io_output_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_output_bits_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_free; // @[ReadMemoryController.scala 251:28]
  ArbiterTree_1 in_arb ( // @[ReadMemoryController.scala 221:25]
    .clock(in_arb_clock),
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_address(in_arb_io_in_0_bits_address),
    .io_in_0_bits_taskID(in_arb_io_in_0_bits_taskID),
    .io_in_1_ready(in_arb_io_in_1_ready),
    .io_in_1_valid(in_arb_io_in_1_valid),
    .io_in_1_bits_address(in_arb_io_in_1_bits_address),
    .io_in_1_bits_taskID(in_arb_io_in_1_bits_taskID),
    .io_in_2_ready(in_arb_io_in_2_ready),
    .io_in_2_valid(in_arb_io_in_2_valid),
    .io_in_2_bits_address(in_arb_io_in_2_bits_address),
    .io_in_2_bits_taskID(in_arb_io_in_2_bits_taskID),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_RouteID(in_arb_io_out_bits_RouteID),
    .io_out_bits_address(in_arb_io_out_bits_address),
    .io_out_bits_taskID(in_arb_io_out_bits_taskID),
    .io_out_bits_Typ(in_arb_io_out_bits_Typ)
  );
  Arbiter alloc_arb ( // @[ReadMemoryController.scala 223:25]
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid)
  );
  Arbiter_1 cachereq_arb ( // @[ReadMemoryController.scala 226:31]
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite)
  );
  Demux cacheresp_demux ( // @[ReadMemoryController.scala 228:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  RRArbiter_1 out_arb ( // @[ReadMemoryController.scala 231:25]
    .clock(out_arb_clock),
    .io_in_0_ready(out_arb_io_in_0_ready),
    .io_in_0_valid(out_arb_io_in_0_valid),
    .io_in_0_bits_RouteID(out_arb_io_in_0_bits_RouteID),
    .io_in_0_bits_data(out_arb_io_in_0_bits_data),
    .io_in_1_ready(out_arb_io_in_1_ready),
    .io_in_1_valid(out_arb_io_in_1_valid),
    .io_in_1_bits_RouteID(out_arb_io_in_1_bits_RouteID),
    .io_in_1_bits_data(out_arb_io_in_1_bits_data),
    .io_out_ready(out_arb_io_out_ready),
    .io_out_valid(out_arb_io_out_valid),
    .io_out_bits_RouteID(out_arb_io_out_bits_RouteID),
    .io_out_bits_data(out_arb_io_out_bits_data),
    .io_chosen(out_arb_io_chosen)
  );
  DeMuxTree_1 out_demux ( // @[ReadMemoryController.scala 232:25]
    .clock(out_demux_clock),
    .reset(out_demux_reset),
    .io_outputs_0_valid(out_demux_io_outputs_0_valid),
    .io_outputs_0_data(out_demux_io_outputs_0_data),
    .io_outputs_1_valid(out_demux_io_outputs_1_valid),
    .io_outputs_1_data(out_demux_io_outputs_1_data),
    .io_outputs_2_valid(out_demux_io_outputs_2_valid),
    .io_outputs_2_data(out_demux_io_outputs_2_data),
    .io_input_RouteID(out_demux_io_input_RouteID),
    .io_input_data(out_demux_io_input_data),
    .io_enable(out_demux_io_enable)
  );
  ReadTableEntry ReadTable_0 ( // @[ReadMemoryController.scala 251:28]
    .clock(ReadTable_0_clock),
    .reset(ReadTable_0_reset),
    .io_NodeReq_ready(ReadTable_0_io_NodeReq_ready),
    .io_NodeReq_valid(ReadTable_0_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(ReadTable_0_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(ReadTable_0_io_NodeReq_bits_address),
    .io_NodeReq_bits_taskID(ReadTable_0_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(ReadTable_0_io_NodeReq_bits_Typ),
    .io_MemReq_ready(ReadTable_0_io_MemReq_ready),
    .io_MemReq_valid(ReadTable_0_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadTable_0_io_MemReq_bits_addr),
    .io_MemReq_bits_tag(ReadTable_0_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadTable_0_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadTable_0_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadTable_0_io_MemResp_valid),
    .io_MemResp_data(ReadTable_0_io_MemResp_data),
    .io_output_ready(ReadTable_0_io_output_ready),
    .io_output_valid(ReadTable_0_io_output_valid),
    .io_output_bits_RouteID(ReadTable_0_io_output_bits_RouteID),
    .io_output_bits_data(ReadTable_0_io_output_bits_data),
    .io_free(ReadTable_0_io_free)
  );
  ReadTableEntry_1 ReadTable_1 ( // @[ReadMemoryController.scala 251:28]
    .clock(ReadTable_1_clock),
    .reset(ReadTable_1_reset),
    .io_NodeReq_ready(ReadTable_1_io_NodeReq_ready),
    .io_NodeReq_valid(ReadTable_1_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(ReadTable_1_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(ReadTable_1_io_NodeReq_bits_address),
    .io_NodeReq_bits_taskID(ReadTable_1_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(ReadTable_1_io_NodeReq_bits_Typ),
    .io_MemReq_ready(ReadTable_1_io_MemReq_ready),
    .io_MemReq_valid(ReadTable_1_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadTable_1_io_MemReq_bits_addr),
    .io_MemReq_bits_tag(ReadTable_1_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadTable_1_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadTable_1_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadTable_1_io_MemResp_valid),
    .io_MemResp_data(ReadTable_1_io_MemResp_data),
    .io_output_ready(ReadTable_1_io_output_ready),
    .io_output_valid(ReadTable_1_io_output_valid),
    .io_output_bits_RouteID(ReadTable_1_io_output_bits_RouteID),
    .io_output_bits_data(ReadTable_1_io_output_bits_data),
    .io_free(ReadTable_1_io_free)
  );
  assign io_ReadIn_0_ready = in_arb_io_in_0_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_1_ready = in_arb_io_in_1_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_2_ready = in_arb_io_in_2_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadOut_0_valid = out_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_0_data = out_demux_io_outputs_0_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_1_valid = out_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_1_data = out_demux_io_outputs_1_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_2_valid = out_demux_io_outputs_2_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_2_data = out_demux_io_outputs_2_data; // @[ReadMemoryController.scala 241:19]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[ReadMemoryController.scala 288:13]
  assign in_arb_clock = clock;
  assign in_arb_io_in_0_valid = io_ReadIn_0_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_0_bits_address = io_ReadIn_0_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_0_bits_taskID = io_ReadIn_0_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_valid = io_ReadIn_1_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_bits_address = io_ReadIn_1_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_bits_taskID = io_ReadIn_1_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_2_valid = io_ReadIn_2_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_2_bits_address = io_ReadIn_2_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_2_bits_taskID = io_ReadIn_2_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_out_ready = alloc_arb_io_out_valid; // @[ReadMemoryController.scala 283:23]
  assign alloc_arb_io_in_0_valid = ReadTable_0_io_free; // @[ReadMemoryController.scala 254:30]
  assign alloc_arb_io_in_1_valid = ReadTable_1_io_free; // @[ReadMemoryController.scala 254:30]
  assign alloc_arb_io_out_ready = in_arb_io_out_valid; // @[ReadMemoryController.scala 284:26]
  assign cachereq_arb_io_in_0_valid = ReadTable_0_io_MemReq_valid; // @[ReadMemoryController.scala 260:33]
  assign cachereq_arb_io_in_0_bits_addr = ReadTable_0_io_MemReq_bits_addr; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_data = 32'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_mask = 4'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_tag = ReadTable_0_io_MemReq_bits_tag; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_taskID = ReadTable_0_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_iswrite = ReadTable_0_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_valid = ReadTable_1_io_MemReq_valid; // @[ReadMemoryController.scala 260:33]
  assign cachereq_arb_io_in_1_bits_addr = ReadTable_1_io_MemReq_bits_addr; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_data = 32'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_mask = 4'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_tag = ReadTable_1_io_MemReq_bits_tag; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_taskID = ReadTable_1_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_iswrite = ReadTable_1_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[ReadMemoryController.scala 288:13]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[ReadMemoryController.scala 291:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[ReadMemoryController.scala 292:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[ReadMemoryController.scala 292:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_tag[0]; // @[ReadMemoryController.scala 293:26]
  assign out_arb_clock = clock;
  assign out_arb_io_in_0_valid = ReadTable_0_io_output_valid; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_0_bits_RouteID = ReadTable_0_io_output_bits_RouteID; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_0_bits_data = ReadTable_0_io_output_bits_data; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_valid = ReadTable_1_io_output_valid; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_bits_RouteID = ReadTable_1_io_output_bits_RouteID; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_bits_data = ReadTable_1_io_output_bits_data; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_out_ready = 1'h1; // @[ReadMemoryController.scala 296:24]
  assign out_demux_clock = clock;
  assign out_demux_reset = reset;
  assign out_demux_io_input_RouteID = out_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 298:22]
  assign out_demux_io_input_data = out_arb_io_out_bits_data; // @[ReadMemoryController.scala 298:22]
  assign out_demux_io_enable = out_arb_io_out_ready & out_arb_io_out_valid; // @[ReadMemoryController.scala 297:23]
  assign ReadTable_0_clock = clock;
  assign ReadTable_0_reset = reset;
  assign ReadTable_0_io_NodeReq_valid = alloc_arb_io_in_0_ready & alloc_arb_io_in_0_valid; // @[ReadMemoryController.scala 256:33]
  assign ReadTable_0_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_MemReq_ready = cachereq_arb_io_in_0_ready; // @[ReadMemoryController.scala 262:32]
  assign ReadTable_0_io_MemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_0_io_MemResp_data = cacheresp_demux_io_outputs_0_data; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_0_io_output_ready = out_arb_io_in_0_ready; // @[ReadMemoryController.scala 268:22]
  assign ReadTable_1_clock = clock;
  assign ReadTable_1_reset = reset;
  assign ReadTable_1_io_NodeReq_valid = alloc_arb_io_in_1_ready & alloc_arb_io_in_1_valid; // @[ReadMemoryController.scala 256:33]
  assign ReadTable_1_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_MemReq_ready = cachereq_arb_io_in_1_ready; // @[ReadMemoryController.scala 262:32]
  assign ReadTable_1_io_MemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_1_io_MemResp_data = cacheresp_demux_io_outputs_1_data; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_1_io_output_ready = out_arb_io_in_1_ready; // @[ReadMemoryController.scala 268:22]
endmodule
module RRArbiter_2(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_data,
  input  [3:0]  io_in_0_bits_mask,
  input  [7:0]  io_in_0_bits_tag,
  input  [9:0]  io_in_0_bits_taskID,
  input         io_in_0_bits_iswrite,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_data,
  input  [3:0]  io_in_1_bits_mask,
  input  [7:0]  io_in_1_bits_tag,
  input  [9:0]  io_in_1_bits_taskID,
  input         io_in_1_bits_iswrite,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_data,
  output [3:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [9:0]  io_out_bits_taskID,
  output        io_out_bits_iswrite,
  output        io_chosen
);
  wire  _T_79; // @[Decoupled.scala 37:37]
  reg  _T_81; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  wire  _T_84; // @[Arbiter.scala 67:57]
  wire  _T_86; // @[Arbiter.scala 68:83]
  wire  _T_89; // @[Arbiter.scala 31:68]
  wire  _T_93; // @[Arbiter.scala 31:78]
  wire  _T_95; // @[Arbiter.scala 31:78]
  wire  _T_99; // @[Arbiter.scala 72:50]
  wire  _GEN_19; // @[Arbiter.scala 77:27]
  assign _T_79 = io_out_ready & io_out_valid; // @[Decoupled.scala 37:37]
  assign _T_84 = 1'h1 > _T_81; // @[Arbiter.scala 67:57]
  assign _T_86 = io_in_1_valid & _T_84; // @[Arbiter.scala 68:83]
  assign _T_89 = _T_86 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_93 = _T_86 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_95 = _T_89 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_99 = _T_84 | _T_95; // @[Arbiter.scala 72:50]
  assign _GEN_19 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_93 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_99 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_mask = io_chosen ? io_in_1_bits_mask : io_in_0_bits_mask; // @[Arbiter.scala 42:15]
  assign io_out_bits_tag = io_chosen ? io_in_1_bits_tag : io_in_0_bits_tag; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_iswrite = io_chosen ? io_in_1_bits_iswrite : io_in_0_bits_iswrite; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_86 ? 1'h1 : _GEN_19; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_81 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_79) begin
      _T_81 <= io_chosen;
    end
  end
endmodule
module ReadWriteArbiter(
  input         clock,
  output        io_ReadMemReq_ready,
  input         io_ReadMemReq_valid,
  input  [31:0] io_ReadMemReq_bits_addr,
  input  [31:0] io_ReadMemReq_bits_data,
  input  [3:0]  io_ReadMemReq_bits_mask,
  input  [7:0]  io_ReadMemReq_bits_tag,
  input  [9:0]  io_ReadMemReq_bits_taskID,
  input         io_ReadMemReq_bits_iswrite,
  output        io_WriteMemReq_ready,
  input         io_WriteMemReq_valid,
  input  [31:0] io_WriteMemReq_bits_addr,
  input  [31:0] io_WriteMemReq_bits_data,
  input  [3:0]  io_WriteMemReq_bits_mask,
  input  [7:0]  io_WriteMemReq_bits_tag,
  input  [9:0]  io_WriteMemReq_bits_taskID,
  input         io_WriteMemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  output        io_ReadMemResp_valid,
  output [31:0] io_ReadMemResp_bits_data,
  output [7:0]  io_ReadMemResp_bits_tag,
  output        io_WriteMemResp_valid,
  output [31:0] io_WriteMemResp_bits_data,
  output [7:0]  io_WriteMemResp_bits_tag,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite
);
  wire  cachereq_arb_clock; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [9:0] cachereq_arb_io_in_0_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [9:0] cachereq_arb_io_in_1_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [9:0] cachereq_arb_io_out_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_chosen; // @[ReadWriteArbiter.scala 48:31]
  wire  cacheresp_demux_io_en; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_sel; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[ReadWriteArbiter.scala 50:31]
  RRArbiter_2 cachereq_arb ( // @[ReadWriteArbiter.scala 48:31]
    .clock(cachereq_arb_clock),
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite),
    .io_chosen(cachereq_arb_io_chosen)
  );
  Demux cacheresp_demux ( // @[ReadWriteArbiter.scala 50:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  assign io_ReadMemReq_ready = cachereq_arb_io_in_0_ready; // @[ReadWriteArbiter.scala 57:29]
  assign io_WriteMemReq_ready = cachereq_arb_io_in_1_ready; // @[ReadWriteArbiter.scala 58:29]
  assign io_ReadMemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[ReadWriteArbiter.scala 69:24]
  assign io_ReadMemResp_bits_data = cacheresp_demux_io_outputs_0_data; // @[ReadWriteArbiter.scala 68:23]
  assign io_ReadMemResp_bits_tag = cacheresp_demux_io_outputs_0_tag; // @[ReadWriteArbiter.scala 68:23]
  assign io_WriteMemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[ReadWriteArbiter.scala 71:25]
  assign io_WriteMemResp_bits_data = cacheresp_demux_io_outputs_1_data; // @[ReadWriteArbiter.scala 70:24]
  assign io_WriteMemResp_bits_tag = cacheresp_demux_io_outputs_1_tag; // @[ReadWriteArbiter.scala 70:24]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[ReadWriteArbiter.scala 62:19]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[ReadWriteArbiter.scala 61:18]
  assign cachereq_arb_clock = clock;
  assign cachereq_arb_io_in_0_valid = io_ReadMemReq_valid; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_addr = io_ReadMemReq_bits_addr; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_data = io_ReadMemReq_bits_data; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_mask = io_ReadMemReq_bits_mask; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_tag = io_ReadMemReq_bits_tag; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_taskID = io_ReadMemReq_bits_taskID; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_iswrite = io_ReadMemReq_bits_iswrite; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_1_valid = io_WriteMemReq_valid; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_addr = io_WriteMemReq_bits_addr; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_data = io_WriteMemReq_bits_data; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_mask = io_WriteMemReq_bits_mask; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_tag = io_WriteMemReq_bits_tag; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_taskID = io_WriteMemReq_bits_taskID; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_iswrite = io_WriteMemReq_bits_iswrite; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[ReadWriteArbiter.scala 60:29]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[ReadWriteArbiter.scala 76:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[ReadWriteArbiter.scala 77:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[ReadWriteArbiter.scala 77:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_iswrite; // @[ReadWriteArbiter.scala 80:26]
endmodule
module UnifiedController(
  input         clock,
  input         reset,
  output        io_WriteIn_0_ready,
  input         io_WriteIn_0_valid,
  input  [21:0] io_WriteIn_0_bits_address,
  input  [31:0] io_WriteIn_0_bits_data,
  input  [9:0]  io_WriteIn_0_bits_taskID,
  output        io_WriteOut_0_valid,
  output        io_ReadIn_0_ready,
  input         io_ReadIn_0_valid,
  input  [31:0] io_ReadIn_0_bits_address,
  input  [9:0]  io_ReadIn_0_bits_taskID,
  output        io_ReadIn_1_ready,
  input         io_ReadIn_1_valid,
  input  [31:0] io_ReadIn_1_bits_address,
  input  [9:0]  io_ReadIn_1_bits_taskID,
  output        io_ReadIn_2_ready,
  input         io_ReadIn_2_valid,
  input  [31:0] io_ReadIn_2_bits_address,
  input  [9:0]  io_ReadIn_2_bits_taskID,
  output        io_ReadOut_0_valid,
  output [31:0] io_ReadOut_0_data,
  output        io_ReadOut_1_valid,
  output [31:0] io_ReadOut_1_data,
  output        io_ReadOut_2_valid,
  output [31:0] io_ReadOut_2_data,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite
);
  wire  WriteController_clock; // @[UnifiedController.scala 64:32]
  wire  WriteController_reset; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_WriteIn_0_ready; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_WriteIn_0_valid; // @[UnifiedController.scala 64:32]
  wire [21:0] WriteController_io_WriteIn_0_bits_address; // @[UnifiedController.scala 64:32]
  wire [31:0] WriteController_io_WriteIn_0_bits_data; // @[UnifiedController.scala 64:32]
  wire [9:0] WriteController_io_WriteIn_0_bits_taskID; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_WriteOut_0_valid; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_MemReq_ready; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_MemReq_valid; // @[UnifiedController.scala 64:32]
  wire [31:0] WriteController_io_MemReq_bits_addr; // @[UnifiedController.scala 64:32]
  wire [31:0] WriteController_io_MemReq_bits_data; // @[UnifiedController.scala 64:32]
  wire [3:0] WriteController_io_MemReq_bits_mask; // @[UnifiedController.scala 64:32]
  wire [7:0] WriteController_io_MemReq_bits_tag; // @[UnifiedController.scala 64:32]
  wire [9:0] WriteController_io_MemReq_bits_taskID; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 64:32]
  wire  WriteController_io_MemResp_valid; // @[UnifiedController.scala 64:32]
  wire [31:0] WriteController_io_MemResp_bits_data; // @[UnifiedController.scala 64:32]
  wire [7:0] WriteController_io_MemResp_bits_tag; // @[UnifiedController.scala 64:32]
  wire  ReadController_clock; // @[UnifiedController.scala 65:32]
  wire  ReadController_reset; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadIn_0_ready; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadIn_0_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_ReadIn_0_bits_address; // @[UnifiedController.scala 65:32]
  wire [9:0] ReadController_io_ReadIn_0_bits_taskID; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadIn_1_ready; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadIn_1_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_ReadIn_1_bits_address; // @[UnifiedController.scala 65:32]
  wire [9:0] ReadController_io_ReadIn_1_bits_taskID; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadIn_2_ready; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadIn_2_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_ReadIn_2_bits_address; // @[UnifiedController.scala 65:32]
  wire [9:0] ReadController_io_ReadIn_2_bits_taskID; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadOut_0_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_ReadOut_0_data; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadOut_1_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_ReadOut_1_data; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_ReadOut_2_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_ReadOut_2_data; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_MemReq_ready; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_MemReq_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_MemReq_bits_addr; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_MemReq_bits_data; // @[UnifiedController.scala 65:32]
  wire [3:0] ReadController_io_MemReq_bits_mask; // @[UnifiedController.scala 65:32]
  wire [7:0] ReadController_io_MemReq_bits_tag; // @[UnifiedController.scala 65:32]
  wire [9:0] ReadController_io_MemReq_bits_taskID; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 65:32]
  wire  ReadController_io_MemResp_valid; // @[UnifiedController.scala 65:32]
  wire [31:0] ReadController_io_MemResp_bits_data; // @[UnifiedController.scala 65:32]
  wire [7:0] ReadController_io_MemResp_bits_tag; // @[UnifiedController.scala 65:32]
  wire  ReadWriteArbiter_clock; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_ReadMemReq_ready; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_ReadMemReq_valid; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemReq_bits_addr; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemReq_bits_data; // @[UnifiedController.scala 66:32]
  wire [3:0] ReadWriteArbiter_io_ReadMemReq_bits_mask; // @[UnifiedController.scala 66:32]
  wire [7:0] ReadWriteArbiter_io_ReadMemReq_bits_tag; // @[UnifiedController.scala 66:32]
  wire [9:0] ReadWriteArbiter_io_ReadMemReq_bits_taskID; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_ReadMemReq_bits_iswrite; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_WriteMemReq_ready; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_WriteMemReq_valid; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemReq_bits_addr; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemReq_bits_data; // @[UnifiedController.scala 66:32]
  wire [3:0] ReadWriteArbiter_io_WriteMemReq_bits_mask; // @[UnifiedController.scala 66:32]
  wire [7:0] ReadWriteArbiter_io_WriteMemReq_bits_tag; // @[UnifiedController.scala 66:32]
  wire [9:0] ReadWriteArbiter_io_WriteMemReq_bits_taskID; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_WriteMemReq_bits_iswrite; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_MemResp_valid; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_MemResp_bits_data; // @[UnifiedController.scala 66:32]
  wire [7:0] ReadWriteArbiter_io_MemResp_bits_tag; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_MemResp_bits_iswrite; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_ReadMemResp_valid; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemResp_bits_data; // @[UnifiedController.scala 66:32]
  wire [7:0] ReadWriteArbiter_io_ReadMemResp_bits_tag; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_WriteMemResp_valid; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemResp_bits_data; // @[UnifiedController.scala 66:32]
  wire [7:0] ReadWriteArbiter_io_WriteMemResp_bits_tag; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_MemReq_ready; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_MemReq_valid; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_MemReq_bits_addr; // @[UnifiedController.scala 66:32]
  wire [31:0] ReadWriteArbiter_io_MemReq_bits_data; // @[UnifiedController.scala 66:32]
  wire [3:0] ReadWriteArbiter_io_MemReq_bits_mask; // @[UnifiedController.scala 66:32]
  wire [7:0] ReadWriteArbiter_io_MemReq_bits_tag; // @[UnifiedController.scala 66:32]
  wire [9:0] ReadWriteArbiter_io_MemReq_bits_taskID; // @[UnifiedController.scala 66:32]
  wire  ReadWriteArbiter_io_MemReq_bits_iswrite; // @[UnifiedController.scala 66:32]
  WriteMemoryController WriteController ( // @[UnifiedController.scala 64:32]
    .clock(WriteController_clock),
    .reset(WriteController_reset),
    .io_WriteIn_0_ready(WriteController_io_WriteIn_0_ready),
    .io_WriteIn_0_valid(WriteController_io_WriteIn_0_valid),
    .io_WriteIn_0_bits_address(WriteController_io_WriteIn_0_bits_address),
    .io_WriteIn_0_bits_data(WriteController_io_WriteIn_0_bits_data),
    .io_WriteIn_0_bits_taskID(WriteController_io_WriteIn_0_bits_taskID),
    .io_WriteOut_0_valid(WriteController_io_WriteOut_0_valid),
    .io_MemReq_ready(WriteController_io_MemReq_ready),
    .io_MemReq_valid(WriteController_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteController_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteController_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteController_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(WriteController_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(WriteController_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteController_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteController_io_MemResp_valid),
    .io_MemResp_bits_data(WriteController_io_MemResp_bits_data),
    .io_MemResp_bits_tag(WriteController_io_MemResp_bits_tag)
  );
  ReadMemoryController ReadController ( // @[UnifiedController.scala 65:32]
    .clock(ReadController_clock),
    .reset(ReadController_reset),
    .io_ReadIn_0_ready(ReadController_io_ReadIn_0_ready),
    .io_ReadIn_0_valid(ReadController_io_ReadIn_0_valid),
    .io_ReadIn_0_bits_address(ReadController_io_ReadIn_0_bits_address),
    .io_ReadIn_0_bits_taskID(ReadController_io_ReadIn_0_bits_taskID),
    .io_ReadIn_1_ready(ReadController_io_ReadIn_1_ready),
    .io_ReadIn_1_valid(ReadController_io_ReadIn_1_valid),
    .io_ReadIn_1_bits_address(ReadController_io_ReadIn_1_bits_address),
    .io_ReadIn_1_bits_taskID(ReadController_io_ReadIn_1_bits_taskID),
    .io_ReadIn_2_ready(ReadController_io_ReadIn_2_ready),
    .io_ReadIn_2_valid(ReadController_io_ReadIn_2_valid),
    .io_ReadIn_2_bits_address(ReadController_io_ReadIn_2_bits_address),
    .io_ReadIn_2_bits_taskID(ReadController_io_ReadIn_2_bits_taskID),
    .io_ReadOut_0_valid(ReadController_io_ReadOut_0_valid),
    .io_ReadOut_0_data(ReadController_io_ReadOut_0_data),
    .io_ReadOut_1_valid(ReadController_io_ReadOut_1_valid),
    .io_ReadOut_1_data(ReadController_io_ReadOut_1_data),
    .io_ReadOut_2_valid(ReadController_io_ReadOut_2_valid),
    .io_ReadOut_2_data(ReadController_io_ReadOut_2_data),
    .io_MemReq_ready(ReadController_io_MemReq_ready),
    .io_MemReq_valid(ReadController_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadController_io_MemReq_bits_addr),
    .io_MemReq_bits_data(ReadController_io_MemReq_bits_data),
    .io_MemReq_bits_mask(ReadController_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(ReadController_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadController_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadController_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadController_io_MemResp_valid),
    .io_MemResp_bits_data(ReadController_io_MemResp_bits_data),
    .io_MemResp_bits_tag(ReadController_io_MemResp_bits_tag)
  );
  ReadWriteArbiter ReadWriteArbiter ( // @[UnifiedController.scala 66:32]
    .clock(ReadWriteArbiter_clock),
    .io_ReadMemReq_ready(ReadWriteArbiter_io_ReadMemReq_ready),
    .io_ReadMemReq_valid(ReadWriteArbiter_io_ReadMemReq_valid),
    .io_ReadMemReq_bits_addr(ReadWriteArbiter_io_ReadMemReq_bits_addr),
    .io_ReadMemReq_bits_data(ReadWriteArbiter_io_ReadMemReq_bits_data),
    .io_ReadMemReq_bits_mask(ReadWriteArbiter_io_ReadMemReq_bits_mask),
    .io_ReadMemReq_bits_tag(ReadWriteArbiter_io_ReadMemReq_bits_tag),
    .io_ReadMemReq_bits_taskID(ReadWriteArbiter_io_ReadMemReq_bits_taskID),
    .io_ReadMemReq_bits_iswrite(ReadWriteArbiter_io_ReadMemReq_bits_iswrite),
    .io_WriteMemReq_ready(ReadWriteArbiter_io_WriteMemReq_ready),
    .io_WriteMemReq_valid(ReadWriteArbiter_io_WriteMemReq_valid),
    .io_WriteMemReq_bits_addr(ReadWriteArbiter_io_WriteMemReq_bits_addr),
    .io_WriteMemReq_bits_data(ReadWriteArbiter_io_WriteMemReq_bits_data),
    .io_WriteMemReq_bits_mask(ReadWriteArbiter_io_WriteMemReq_bits_mask),
    .io_WriteMemReq_bits_tag(ReadWriteArbiter_io_WriteMemReq_bits_tag),
    .io_WriteMemReq_bits_taskID(ReadWriteArbiter_io_WriteMemReq_bits_taskID),
    .io_WriteMemReq_bits_iswrite(ReadWriteArbiter_io_WriteMemReq_bits_iswrite),
    .io_MemResp_valid(ReadWriteArbiter_io_MemResp_valid),
    .io_MemResp_bits_data(ReadWriteArbiter_io_MemResp_bits_data),
    .io_MemResp_bits_tag(ReadWriteArbiter_io_MemResp_bits_tag),
    .io_MemResp_bits_iswrite(ReadWriteArbiter_io_MemResp_bits_iswrite),
    .io_ReadMemResp_valid(ReadWriteArbiter_io_ReadMemResp_valid),
    .io_ReadMemResp_bits_data(ReadWriteArbiter_io_ReadMemResp_bits_data),
    .io_ReadMemResp_bits_tag(ReadWriteArbiter_io_ReadMemResp_bits_tag),
    .io_WriteMemResp_valid(ReadWriteArbiter_io_WriteMemResp_valid),
    .io_WriteMemResp_bits_data(ReadWriteArbiter_io_WriteMemResp_bits_data),
    .io_WriteMemResp_bits_tag(ReadWriteArbiter_io_WriteMemResp_bits_tag),
    .io_MemReq_ready(ReadWriteArbiter_io_MemReq_ready),
    .io_MemReq_valid(ReadWriteArbiter_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadWriteArbiter_io_MemReq_bits_addr),
    .io_MemReq_bits_data(ReadWriteArbiter_io_MemReq_bits_data),
    .io_MemReq_bits_mask(ReadWriteArbiter_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(ReadWriteArbiter_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadWriteArbiter_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadWriteArbiter_io_MemReq_bits_iswrite)
  );
  assign io_WriteIn_0_ready = WriteController_io_WriteIn_0_ready; // @[UnifiedController.scala 74:35]
  assign io_WriteOut_0_valid = WriteController_io_WriteOut_0_valid; // @[UnifiedController.scala 75:20]
  assign io_ReadIn_0_ready = ReadController_io_ReadIn_0_ready; // @[UnifiedController.scala 80:33]
  assign io_ReadIn_1_ready = ReadController_io_ReadIn_1_ready; // @[UnifiedController.scala 80:33]
  assign io_ReadIn_2_ready = ReadController_io_ReadIn_2_ready; // @[UnifiedController.scala 80:33]
  assign io_ReadOut_0_valid = ReadController_io_ReadOut_0_valid; // @[UnifiedController.scala 81:19]
  assign io_ReadOut_0_data = ReadController_io_ReadOut_0_data; // @[UnifiedController.scala 81:19]
  assign io_ReadOut_1_valid = ReadController_io_ReadOut_1_valid; // @[UnifiedController.scala 81:19]
  assign io_ReadOut_1_data = ReadController_io_ReadOut_1_data; // @[UnifiedController.scala 81:19]
  assign io_ReadOut_2_valid = ReadController_io_ReadOut_2_valid; // @[UnifiedController.scala 81:19]
  assign io_ReadOut_2_data = ReadController_io_ReadOut_2_data; // @[UnifiedController.scala 81:19]
  assign io_MemReq_valid = ReadWriteArbiter_io_MemReq_valid; // @[UnifiedController.scala 94:19]
  assign io_MemReq_bits_addr = ReadWriteArbiter_io_MemReq_bits_addr; // @[UnifiedController.scala 93:18]
  assign io_MemReq_bits_data = ReadWriteArbiter_io_MemReq_bits_data; // @[UnifiedController.scala 93:18]
  assign io_MemReq_bits_mask = ReadWriteArbiter_io_MemReq_bits_mask; // @[UnifiedController.scala 93:18]
  assign io_MemReq_bits_tag = ReadWriteArbiter_io_MemReq_bits_tag; // @[UnifiedController.scala 93:18]
  assign io_MemReq_bits_taskID = ReadWriteArbiter_io_MemReq_bits_taskID; // @[UnifiedController.scala 93:18]
  assign io_MemReq_bits_iswrite = ReadWriteArbiter_io_MemReq_bits_iswrite; // @[UnifiedController.scala 93:18]
  assign WriteController_clock = clock;
  assign WriteController_reset = reset;
  assign WriteController_io_WriteIn_0_valid = io_WriteIn_0_valid; // @[UnifiedController.scala 74:35]
  assign WriteController_io_WriteIn_0_bits_address = io_WriteIn_0_bits_address; // @[UnifiedController.scala 74:35]
  assign WriteController_io_WriteIn_0_bits_data = io_WriteIn_0_bits_data; // @[UnifiedController.scala 74:35]
  assign WriteController_io_WriteIn_0_bits_taskID = io_WriteIn_0_bits_taskID; // @[UnifiedController.scala 74:35]
  assign WriteController_io_MemReq_ready = ReadWriteArbiter_io_WriteMemReq_ready; // @[UnifiedController.scala 88:35]
  assign WriteController_io_MemResp_valid = ReadWriteArbiter_io_WriteMemResp_valid; // @[UnifiedController.scala 89:30]
  assign WriteController_io_MemResp_bits_data = ReadWriteArbiter_io_WriteMemResp_bits_data; // @[UnifiedController.scala 89:30]
  assign WriteController_io_MemResp_bits_tag = ReadWriteArbiter_io_WriteMemResp_bits_tag; // @[UnifiedController.scala 89:30]
  assign ReadController_clock = clock;
  assign ReadController_reset = reset;
  assign ReadController_io_ReadIn_0_valid = io_ReadIn_0_valid; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_0_bits_address = io_ReadIn_0_bits_address; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_0_bits_taskID = io_ReadIn_0_bits_taskID; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_1_valid = io_ReadIn_1_valid; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_1_bits_address = io_ReadIn_1_bits_address; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_1_bits_taskID = io_ReadIn_1_bits_taskID; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_2_valid = io_ReadIn_2_valid; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_2_bits_address = io_ReadIn_2_bits_address; // @[UnifiedController.scala 80:33]
  assign ReadController_io_ReadIn_2_bits_taskID = io_ReadIn_2_bits_taskID; // @[UnifiedController.scala 80:33]
  assign ReadController_io_MemReq_ready = ReadWriteArbiter_io_ReadMemReq_ready; // @[UnifiedController.scala 85:34]
  assign ReadController_io_MemResp_valid = ReadWriteArbiter_io_ReadMemResp_valid; // @[UnifiedController.scala 86:29]
  assign ReadController_io_MemResp_bits_data = ReadWriteArbiter_io_ReadMemResp_bits_data; // @[UnifiedController.scala 86:29]
  assign ReadController_io_MemResp_bits_tag = ReadWriteArbiter_io_ReadMemResp_bits_tag; // @[UnifiedController.scala 86:29]
  assign ReadWriteArbiter_clock = clock;
  assign ReadWriteArbiter_io_ReadMemReq_valid = ReadController_io_MemReq_valid; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_addr = ReadController_io_MemReq_bits_addr; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_data = ReadController_io_MemReq_bits_data; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_mask = ReadController_io_MemReq_bits_mask; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_tag = ReadController_io_MemReq_bits_tag; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_taskID = ReadController_io_MemReq_bits_taskID; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_iswrite = ReadController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 85:34]
  assign ReadWriteArbiter_io_WriteMemReq_valid = WriteController_io_MemReq_valid; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_addr = WriteController_io_MemReq_bits_addr; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_data = WriteController_io_MemReq_bits_data; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_mask = WriteController_io_MemReq_bits_mask; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_tag = WriteController_io_MemReq_bits_tag; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_taskID = WriteController_io_MemReq_bits_taskID; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_iswrite = WriteController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 88:35]
  assign ReadWriteArbiter_io_MemResp_valid = io_MemResp_valid; // @[UnifiedController.scala 95:31]
  assign ReadWriteArbiter_io_MemResp_bits_data = io_MemResp_bits_data; // @[UnifiedController.scala 95:31]
  assign ReadWriteArbiter_io_MemResp_bits_tag = io_MemResp_bits_tag; // @[UnifiedController.scala 95:31]
  assign ReadWriteArbiter_io_MemResp_bits_iswrite = io_MemResp_bits_iswrite; // @[UnifiedController.scala 95:31]
  assign ReadWriteArbiter_io_MemReq_ready = io_MemReq_ready; // @[UnifiedController.scala 92:36]
endmodule
module SplitCallNew(
  input         clock,
  input         reset,
  output        io_In_ready,
  input         io_In_valid,
  input  [9:0]  io_In_bits_enable_taskID,
  input         io_In_bits_enable_control,
  input  [9:0]  io_In_bits_data_field2_taskID,
  input  [31:0] io_In_bits_data_field2_data,
  input  [9:0]  io_In_bits_data_field1_taskID,
  input  [31:0] io_In_bits_data_field1_data,
  input  [9:0]  io_In_bits_data_field0_taskID,
  input  [31:0] io_In_bits_data_field0_data,
  input         io_Out_enable_ready,
  output        io_Out_enable_valid,
  output [9:0]  io_Out_enable_bits_taskID,
  output        io_Out_enable_bits_control,
  input         io_Out_data_field2_0_ready,
  output        io_Out_data_field2_0_valid,
  output [9:0]  io_Out_data_field2_0_bits_taskID,
  output [31:0] io_Out_data_field2_0_bits_data,
  input         io_Out_data_field1_0_ready,
  output        io_Out_data_field1_0_valid,
  output [9:0]  io_Out_data_field1_0_bits_taskID,
  output [31:0] io_Out_data_field1_0_bits_data,
  input         io_Out_data_field0_0_ready,
  output        io_Out_data_field0_0_valid,
  output [9:0]  io_Out_data_field0_0_bits_taskID,
  output [31:0] io_Out_data_field0_0_bits_data
);
  reg [9:0] inputReg_enable_taskID; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_0;
  reg  inputReg_enable_control; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_1;
  reg [9:0] inputReg_data_field2_taskID; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_2;
  reg [31:0] inputReg_data_field2_data; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_3;
  reg [9:0] inputReg_data_field1_taskID; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_4;
  reg [31:0] inputReg_data_field1_data; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_5;
  reg [9:0] inputReg_data_field0_taskID; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_6;
  reg [31:0] inputReg_data_field0_data; // @[SplitDecoupled.scala 150:26]
  reg [31:0] _RAND_7;
  reg  enableValidReg; // @[SplitDecoupled.scala 152:31]
  reg [31:0] _RAND_8;
  reg  allValid_0; // @[SplitDecoupled.scala 155:49]
  reg [31:0] _RAND_9;
  reg  allValid_1; // @[SplitDecoupled.scala 155:49]
  reg [31:0] _RAND_10;
  reg  allValid_2; // @[SplitDecoupled.scala 155:49]
  reg [31:0] _RAND_11;
  reg  state; // @[SplitDecoupled.scala 164:22]
  reg [31:0] _RAND_12;
  wire  _T_125; // @[SplitDecoupled.scala 166:24]
  wire  _T_126; // @[Conditional.scala 37:30]
  wire  _T_127; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[SplitDecoupled.scala 170:27]
  wire [9:0] _GEN_1; // @[SplitDecoupled.scala 170:27]
  wire  _GEN_2; // @[SplitDecoupled.scala 170:27]
  wire [9:0] _GEN_4; // @[SplitDecoupled.scala 170:27]
  wire [31:0] _GEN_5; // @[SplitDecoupled.scala 170:27]
  wire [9:0] _GEN_7; // @[SplitDecoupled.scala 170:27]
  wire [31:0] _GEN_8; // @[SplitDecoupled.scala 170:27]
  wire [9:0] _GEN_10; // @[SplitDecoupled.scala 170:27]
  wire [31:0] _GEN_11; // @[SplitDecoupled.scala 170:27]
  wire  _T_129; // @[SplitDecoupled.scala 176:36]
  wire  _T_130; // @[SplitDecoupled.scala 176:36]
  wire  _T_132; // @[SplitDecoupled.scala 176:13]
  wire  _T_134; // @[SplitDecoupled.scala 176:45]
  wire  _T_135; // @[SplitDecoupled.scala 176:42]
  wire  _GEN_12; // @[SplitDecoupled.scala 176:62]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_14; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_15; // @[Conditional.scala 40:58]
  wire  _GEN_16; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_18; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_19; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_21; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_22; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_24; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_25; // @[Conditional.scala 40:58]
  wire  _T_137; // @[SplitDecoupled.scala 184:24]
  wire  _GEN_26; // @[SplitDecoupled.scala 184:45]
  wire  _T_140; // @[SplitDecoupled.scala 187:32]
  wire  _GEN_27; // @[SplitDecoupled.scala 187:69]
  wire  _GEN_28; // @[SplitDecoupled.scala 184:45]
  wire  _T_146; // @[SplitDecoupled.scala 187:32]
  wire  _GEN_29; // @[SplitDecoupled.scala 187:69]
  wire  _GEN_30; // @[SplitDecoupled.scala 184:45]
  wire  _T_152; // @[SplitDecoupled.scala 187:32]
  wire  _GEN_31; // @[SplitDecoupled.scala 187:69]
  wire  _GEN_32; // @[SplitDecoupled.scala 195:41]
  wire  _T_158; // @[SplitDecoupled.scala 198:28]
  wire  _GEN_33; // @[SplitDecoupled.scala 198:51]
  assign _T_125 = state == 1'h0; // @[SplitDecoupled.scala 166:24]
  assign _T_126 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_127 = io_In_ready & io_In_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_127 ? 1'h1 : state; // @[SplitDecoupled.scala 170:27]
  assign _GEN_1 = _T_127 ? io_In_bits_enable_taskID : inputReg_enable_taskID; // @[SplitDecoupled.scala 170:27]
  assign _GEN_2 = _T_127 ? io_In_bits_enable_control : inputReg_enable_control; // @[SplitDecoupled.scala 170:27]
  assign _GEN_4 = _T_127 ? io_In_bits_data_field2_taskID : inputReg_data_field2_taskID; // @[SplitDecoupled.scala 170:27]
  assign _GEN_5 = _T_127 ? io_In_bits_data_field2_data : inputReg_data_field2_data; // @[SplitDecoupled.scala 170:27]
  assign _GEN_7 = _T_127 ? io_In_bits_data_field1_taskID : inputReg_data_field1_taskID; // @[SplitDecoupled.scala 170:27]
  assign _GEN_8 = _T_127 ? io_In_bits_data_field1_data : inputReg_data_field1_data; // @[SplitDecoupled.scala 170:27]
  assign _GEN_10 = _T_127 ? io_In_bits_data_field0_taskID : inputReg_data_field0_taskID; // @[SplitDecoupled.scala 170:27]
  assign _GEN_11 = _T_127 ? io_In_bits_data_field0_data : inputReg_data_field0_data; // @[SplitDecoupled.scala 170:27]
  assign _T_129 = allValid_0 | allValid_1; // @[SplitDecoupled.scala 176:36]
  assign _T_130 = _T_129 | allValid_2; // @[SplitDecoupled.scala 176:36]
  assign _T_132 = _T_130 == 1'h0; // @[SplitDecoupled.scala 176:13]
  assign _T_134 = enableValidReg == 1'h0; // @[SplitDecoupled.scala 176:45]
  assign _T_135 = _T_132 & _T_134; // @[SplitDecoupled.scala 176:42]
  assign _GEN_12 = _T_135 ? 1'h0 : state; // @[SplitDecoupled.scala 176:62]
  assign _GEN_13 = state ? _GEN_12 : state; // @[Conditional.scala 39:67]
  assign _GEN_14 = _T_126 ? _GEN_0 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_15 = _T_126 ? _GEN_1 : inputReg_enable_taskID; // @[Conditional.scala 40:58]
  assign _GEN_16 = _T_126 ? _GEN_2 : inputReg_enable_control; // @[Conditional.scala 40:58]
  assign _GEN_18 = _T_126 ? _GEN_4 : inputReg_data_field2_taskID; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_126 ? _GEN_5 : inputReg_data_field2_data; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_126 ? _GEN_7 : inputReg_data_field1_taskID; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_126 ? _GEN_8 : inputReg_data_field1_data; // @[Conditional.scala 40:58]
  assign _GEN_24 = _T_126 ? _GEN_10 : inputReg_data_field0_taskID; // @[Conditional.scala 40:58]
  assign _GEN_25 = _T_126 ? _GEN_11 : inputReg_data_field0_data; // @[Conditional.scala 40:58]
  assign _T_137 = io_In_valid & _T_125; // @[SplitDecoupled.scala 184:24]
  assign _GEN_26 = _T_137 ? 1'h1 : allValid_0; // @[SplitDecoupled.scala 184:45]
  assign _T_140 = state & io_Out_data_field0_0_ready; // @[SplitDecoupled.scala 187:32]
  assign _GEN_27 = _T_140 ? 1'h0 : _GEN_26; // @[SplitDecoupled.scala 187:69]
  assign _GEN_28 = _T_137 ? 1'h1 : allValid_1; // @[SplitDecoupled.scala 184:45]
  assign _T_146 = state & io_Out_data_field1_0_ready; // @[SplitDecoupled.scala 187:32]
  assign _GEN_29 = _T_146 ? 1'h0 : _GEN_28; // @[SplitDecoupled.scala 187:69]
  assign _GEN_30 = _T_137 ? 1'h1 : allValid_2; // @[SplitDecoupled.scala 184:45]
  assign _T_152 = state & io_Out_data_field2_0_ready; // @[SplitDecoupled.scala 187:32]
  assign _GEN_31 = _T_152 ? 1'h0 : _GEN_30; // @[SplitDecoupled.scala 187:69]
  assign _GEN_32 = _T_137 ? 1'h1 : enableValidReg; // @[SplitDecoupled.scala 195:41]
  assign _T_158 = state & io_Out_enable_ready; // @[SplitDecoupled.scala 198:28]
  assign _GEN_33 = _T_158 ? 1'h0 : _GEN_32; // @[SplitDecoupled.scala 198:51]
  assign io_In_ready = state == 1'h0; // @[SplitDecoupled.scala 166:15]
  assign io_Out_enable_valid = enableValidReg; // @[SplitDecoupled.scala 201:23]
  assign io_Out_enable_bits_taskID = inputReg_enable_taskID; // @[SplitDecoupled.scala 202:22]
  assign io_Out_enable_bits_control = inputReg_enable_control; // @[SplitDecoupled.scala 202:22]
  assign io_Out_data_field2_0_valid = allValid_2; // @[SplitDecoupled.scala 190:40]
  assign io_Out_data_field2_0_bits_taskID = inputReg_data_field2_taskID; // @[SplitDecoupled.scala 191:39]
  assign io_Out_data_field2_0_bits_data = inputReg_data_field2_data; // @[SplitDecoupled.scala 191:39]
  assign io_Out_data_field1_0_valid = allValid_1; // @[SplitDecoupled.scala 190:40]
  assign io_Out_data_field1_0_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 191:39]
  assign io_Out_data_field1_0_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 191:39]
  assign io_Out_data_field0_0_valid = allValid_0; // @[SplitDecoupled.scala 190:40]
  assign io_Out_data_field0_0_bits_taskID = inputReg_data_field0_taskID; // @[SplitDecoupled.scala 191:39]
  assign io_Out_data_field0_0_bits_data = inputReg_data_field0_data; // @[SplitDecoupled.scala 191:39]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inputReg_enable_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inputReg_enable_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inputReg_data_field2_taskID = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inputReg_data_field2_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inputReg_data_field1_taskID = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  inputReg_data_field1_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  inputReg_data_field0_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inputReg_data_field0_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enableValidReg = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  allValid_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  allValid_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  allValid_2 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      inputReg_enable_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_enable_taskID <= io_In_bits_enable_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_enable_control <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_enable_control <= io_In_bits_enable_control;
        end
      end
    end
    if (reset) begin
      inputReg_data_field2_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_data_field2_taskID <= io_In_bits_data_field2_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field2_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_data_field2_data <= io_In_bits_data_field2_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_data_field1_taskID <= io_In_bits_data_field1_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_data_field1_data <= io_In_bits_data_field1_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field0_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_data_field0_taskID <= io_In_bits_data_field0_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field0_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          inputReg_data_field0_data <= io_In_bits_data_field0_data;
        end
      end
    end
    if (reset) begin
      enableValidReg <= 1'h0;
    end else begin
      if (_T_158) begin
        enableValidReg <= 1'h0;
      end else begin
        if (_T_137) begin
          enableValidReg <= 1'h1;
        end
      end
    end
    if (reset) begin
      allValid_0 <= 1'h0;
    end else begin
      if (_T_140) begin
        allValid_0 <= 1'h0;
      end else begin
        if (_T_137) begin
          allValid_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allValid_1 <= 1'h0;
    end else begin
      if (_T_146) begin
        allValid_1 <= 1'h0;
      end else begin
        if (_T_137) begin
          allValid_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allValid_2 <= 1'h0;
    end else begin
      if (_T_152) begin
        allValid_2 <= 1'h0;
      end else begin
        if (_T_137) begin
          allValid_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_127) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_135) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [9:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [9:0]  io_InLiveIn_3_bits_taskID,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [9:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [31:0] io_InLiveIn_5_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field5_1_ready,
  output        io_OutLiveIn_field5_1_valid,
  output [31:0] io_OutLiveIn_field5_1_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [9:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [9:0]  io_OutLiveIn_field3_0_bits_taskID,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [9:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [9:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [9:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [9:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [9:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [9:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [9:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_2;
  reg [9:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_3;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_5;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_6;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_7;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_8;
  reg [9:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [9:0] in_live_in_R_3_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [9:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_17;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_18;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_19;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_20;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_21;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_22;
  reg [9:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_23;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_24;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_25;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_26;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_29;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_30;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_31;
  reg  out_live_in_valid_R_5_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_32;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_33;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_34;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_35;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_36;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_37;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_38;
  reg  out_live_in_fire_R_5_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_39;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_40;
  reg [9:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_41;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_42;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_43;
  reg [9:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_44;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_45;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_46;
  reg [9:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_47;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_48;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_49;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_50;
  wire  _T_653; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[LoopBlock.scala 596:26]
  wire  _GEN_2; // @[LoopBlock.scala 596:26]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_656; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_4; // @[LoopBlock.scala 603:33]
  wire  _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_659; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_662; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[LoopBlock.scala 623:33]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_665; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_15; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_16; // @[LoopBlock.scala 623:33]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_668; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_20; // @[LoopBlock.scala 623:33]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_671; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_23; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_24; // @[LoopBlock.scala 623:33]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_674; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_27; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_28; // @[LoopBlock.scala 623:33]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_677; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_32; // @[LoopBlock.scala 623:33]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_680; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_35; // @[LoopBlock.scala 641:37]
  wire [31:0] _GEN_36; // @[LoopBlock.scala 641:37]
  wire  _GEN_37; // @[LoopBlock.scala 641:37]
  wire  _T_682; // @[Decoupled.scala 37:37]
  wire  _GEN_38; // @[LoopBlock.scala 704:39]
  wire  _T_684; // @[Decoupled.scala 37:37]
  wire  _GEN_39; // @[LoopBlock.scala 708:38]
  wire  _T_686; // @[Decoupled.scala 37:37]
  wire  _GEN_40; // @[LoopBlock.scala 713:33]
  wire  _GEN_41; // @[LoopBlock.scala 713:33]
  wire  _T_689; // @[Decoupled.scala 37:37]
  wire  _GEN_42; // @[LoopBlock.scala 722:57]
  wire  _GEN_43; // @[LoopBlock.scala 722:57]
  wire  _T_692; // @[Decoupled.scala 37:37]
  wire  _GEN_44; // @[LoopBlock.scala 722:57]
  wire  _GEN_45; // @[LoopBlock.scala 722:57]
  wire  _T_695; // @[Decoupled.scala 37:37]
  wire  _GEN_46; // @[LoopBlock.scala 722:57]
  wire  _GEN_47; // @[LoopBlock.scala 722:57]
  wire  _T_698; // @[Decoupled.scala 37:37]
  wire  _GEN_48; // @[LoopBlock.scala 722:57]
  wire  _GEN_49; // @[LoopBlock.scala 722:57]
  wire  _T_701; // @[Decoupled.scala 37:37]
  wire  _GEN_50; // @[LoopBlock.scala 722:57]
  wire  _GEN_51; // @[LoopBlock.scala 722:57]
  wire  _T_704; // @[Decoupled.scala 37:37]
  wire  _GEN_52; // @[LoopBlock.scala 722:57]
  wire  _GEN_53; // @[LoopBlock.scala 722:57]
  wire  _T_707; // @[Decoupled.scala 37:37]
  wire  _GEN_54; // @[LoopBlock.scala 722:57]
  wire  _GEN_55; // @[LoopBlock.scala 722:57]
  wire  _T_710; // @[Decoupled.scala 37:37]
  wire  _GEN_56; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_51;
  wire  _T_714; // @[Conditional.scala 37:30]
  wire  _T_715; // @[LoopBlock.scala 765:35]
  wire  _T_716; // @[LoopBlock.scala 765:35]
  wire  _T_717; // @[LoopBlock.scala 765:35]
  wire  _T_718; // @[LoopBlock.scala 765:35]
  wire  _T_719; // @[LoopBlock.scala 765:35]
  wire  _T_720; // @[LoopBlock.scala 869:28]
  wire  _GEN_58; // @[LoopBlock.scala 870:26]
  wire  _GEN_59; // @[LoopBlock.scala 870:26]
  wire  _GEN_60; // @[LoopBlock.scala 870:26]
  wire  _GEN_61; // @[LoopBlock.scala 870:26]
  wire  _GEN_62; // @[LoopBlock.scala 870:26]
  wire  _GEN_63; // @[LoopBlock.scala 870:26]
  wire  _GEN_64; // @[LoopBlock.scala 870:26]
  wire  _GEN_65; // @[LoopBlock.scala 870:26]
  wire  _GEN_66; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_67; // @[LoopBlock.scala 870:26]
  wire  _GEN_68; // @[LoopBlock.scala 870:26]
  wire  _GEN_69; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_70; // @[LoopBlock.scala 870:26]
  wire  _GEN_71; // @[LoopBlock.scala 870:26]
  wire [1:0] _GEN_72; // @[LoopBlock.scala 870:26]
  wire  _GEN_73; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_74; // @[LoopBlock.scala 870:26]
  wire  _GEN_75; // @[LoopBlock.scala 870:26]
  wire  _GEN_76; // @[LoopBlock.scala 869:48]
  wire  _GEN_77; // @[LoopBlock.scala 869:48]
  wire  _GEN_78; // @[LoopBlock.scala 869:48]
  wire  _GEN_79; // @[LoopBlock.scala 869:48]
  wire  _GEN_80; // @[LoopBlock.scala 869:48]
  wire  _GEN_81; // @[LoopBlock.scala 869:48]
  wire  _GEN_82; // @[LoopBlock.scala 869:48]
  wire  _GEN_83; // @[LoopBlock.scala 869:48]
  wire  _GEN_84; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_85; // @[LoopBlock.scala 869:48]
  wire  _GEN_86; // @[LoopBlock.scala 869:48]
  wire  _GEN_87; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_88; // @[LoopBlock.scala 869:48]
  wire  _GEN_89; // @[LoopBlock.scala 869:48]
  wire [1:0] _GEN_90; // @[LoopBlock.scala 869:48]
  wire  _GEN_91; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_92; // @[LoopBlock.scala 869:48]
  wire  _GEN_93; // @[LoopBlock.scala 869:48]
  wire  _T_742; // @[Conditional.scala 37:30]
  wire  _T_743; // @[LoopBlock.scala 898:30]
  wire  _T_746; // @[LoopBlock.scala 825:65]
  wire  _T_747; // @[LoopBlock.scala 828:26]
  wire  _T_748; // @[LoopBlock.scala 828:26]
  wire  _T_749; // @[LoopBlock.scala 828:26]
  wire  _T_750; // @[LoopBlock.scala 828:26]
  wire  _T_751; // @[LoopBlock.scala 828:26]
  wire  _T_752; // @[LoopBlock.scala 899:29]
  wire  _GEN_94; // @[LoopBlock.scala 936:64]
  wire  _GEN_95; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_96; // @[LoopBlock.scala 936:64]
  wire  _GEN_97; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_98; // @[LoopBlock.scala 936:64]
  wire  _GEN_99; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_100; // @[LoopBlock.scala 936:64]
  wire [1:0] _GEN_101; // @[LoopBlock.scala 936:64]
  wire  _GEN_102; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_103; // @[LoopBlock.scala 903:56]
  wire  _GEN_104; // @[LoopBlock.scala 903:56]
  wire  _GEN_105; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_106; // @[LoopBlock.scala 903:56]
  wire  _GEN_107; // @[LoopBlock.scala 903:56]
  wire  _GEN_108; // @[LoopBlock.scala 903:56]
  wire  _GEN_109; // @[LoopBlock.scala 903:56]
  wire  _GEN_110; // @[LoopBlock.scala 903:56]
  wire  _GEN_111; // @[LoopBlock.scala 903:56]
  wire  _GEN_112; // @[LoopBlock.scala 903:56]
  wire  _GEN_113; // @[LoopBlock.scala 903:56]
  wire  _GEN_114; // @[LoopBlock.scala 903:56]
  wire  _GEN_116; // @[LoopBlock.scala 903:56]
  wire  _GEN_117; // @[LoopBlock.scala 903:56]
  wire  _GEN_118; // @[LoopBlock.scala 903:56]
  wire  _GEN_119; // @[LoopBlock.scala 903:56]
  wire  _GEN_120; // @[LoopBlock.scala 903:56]
  wire  _GEN_121; // @[LoopBlock.scala 903:56]
  wire  _GEN_122; // @[LoopBlock.scala 903:56]
  wire  _GEN_123; // @[LoopBlock.scala 903:56]
  wire  _GEN_124; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_125; // @[LoopBlock.scala 903:56]
  wire  _GEN_126; // @[LoopBlock.scala 903:56]
  wire  _GEN_127; // @[LoopBlock.scala 903:56]
  wire  _GEN_129; // @[LoopBlock.scala 903:56]
  wire  _GEN_130; // @[LoopBlock.scala 903:56]
  wire [1:0] _GEN_131; // @[LoopBlock.scala 903:56]
  wire  _GEN_132; // @[LoopBlock.scala 903:56]
  wire  _GEN_133; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_134; // @[LoopBlock.scala 903:56]
  wire  _GEN_135; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_136; // @[LoopBlock.scala 900:55]
  wire  _GEN_137; // @[LoopBlock.scala 900:55]
  wire  _GEN_138; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_139; // @[LoopBlock.scala 900:55]
  wire  _GEN_140; // @[LoopBlock.scala 900:55]
  wire  _GEN_141; // @[LoopBlock.scala 900:55]
  wire  _GEN_142; // @[LoopBlock.scala 900:55]
  wire  _GEN_143; // @[LoopBlock.scala 900:55]
  wire  _GEN_144; // @[LoopBlock.scala 900:55]
  wire  _GEN_145; // @[LoopBlock.scala 900:55]
  wire  _GEN_146; // @[LoopBlock.scala 900:55]
  wire  _GEN_147; // @[LoopBlock.scala 900:55]
  wire  _GEN_149; // @[LoopBlock.scala 900:55]
  wire  _GEN_150; // @[LoopBlock.scala 900:55]
  wire  _GEN_151; // @[LoopBlock.scala 900:55]
  wire  _GEN_152; // @[LoopBlock.scala 900:55]
  wire  _GEN_153; // @[LoopBlock.scala 900:55]
  wire  _GEN_154; // @[LoopBlock.scala 900:55]
  wire  _GEN_155; // @[LoopBlock.scala 900:55]
  wire  _GEN_156; // @[LoopBlock.scala 900:55]
  wire  _GEN_157; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_158; // @[LoopBlock.scala 900:55]
  wire  _GEN_159; // @[LoopBlock.scala 900:55]
  wire  _GEN_160; // @[LoopBlock.scala 900:55]
  wire  _GEN_162; // @[LoopBlock.scala 900:55]
  wire  _GEN_163; // @[LoopBlock.scala 900:55]
  wire [1:0] _GEN_164; // @[LoopBlock.scala 900:55]
  wire  _GEN_165; // @[LoopBlock.scala 900:55]
  wire  _GEN_166; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_167; // @[LoopBlock.scala 900:55]
  wire  _T_805; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_168; // @[LoopBlock.scala 955:48]
  wire  _GEN_169; // @[LoopBlock.scala 955:48]
  wire  _GEN_170; // @[LoopBlock.scala 955:48]
  wire  _GEN_171; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_172; // @[LoopBlock.scala 955:48]
  wire  _GEN_173; // @[LoopBlock.scala 955:48]
  wire  _GEN_174; // @[LoopBlock.scala 955:48]
  wire  _GEN_176; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_177; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_180; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_181; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_183; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_186; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_187; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_189; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_190; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_192; // @[LoopBlock.scala 955:48]
  wire  _GEN_195; // @[LoopBlock.scala 955:48]
  wire  _GEN_196; // @[LoopBlock.scala 955:48]
  wire  _GEN_197; // @[LoopBlock.scala 955:48]
  wire  _GEN_198; // @[LoopBlock.scala 955:48]
  wire  _GEN_199; // @[LoopBlock.scala 955:48]
  wire  _GEN_200; // @[LoopBlock.scala 955:48]
  wire  _GEN_201; // @[LoopBlock.scala 955:48]
  wire [1:0] _GEN_202; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_203; // @[Conditional.scala 39:67]
  wire  _GEN_204; // @[Conditional.scala 39:67]
  wire  _GEN_205; // @[Conditional.scala 39:67]
  wire  _GEN_206; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_207; // @[Conditional.scala 39:67]
  wire  _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_209; // @[Conditional.scala 39:67]
  wire  _GEN_211; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_212; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_215; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_216; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_218; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_221; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_222; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_224; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_225; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_227; // @[Conditional.scala 39:67]
  wire  _GEN_230; // @[Conditional.scala 39:67]
  wire  _GEN_231; // @[Conditional.scala 39:67]
  wire  _GEN_232; // @[Conditional.scala 39:67]
  wire  _GEN_233; // @[Conditional.scala 39:67]
  wire  _GEN_234; // @[Conditional.scala 39:67]
  wire  _GEN_235; // @[Conditional.scala 39:67]
  wire  _GEN_236; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_237; // @[Conditional.scala 39:67]
  wire  _GEN_238; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_239; // @[Conditional.scala 39:67]
  wire  _GEN_240; // @[Conditional.scala 39:67]
  wire  _GEN_241; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_242; // @[Conditional.scala 39:67]
  wire  _GEN_243; // @[Conditional.scala 39:67]
  wire  _GEN_244; // @[Conditional.scala 39:67]
  wire  _GEN_245; // @[Conditional.scala 39:67]
  wire  _GEN_246; // @[Conditional.scala 39:67]
  wire  _GEN_247; // @[Conditional.scala 39:67]
  wire  _GEN_248; // @[Conditional.scala 39:67]
  wire  _GEN_249; // @[Conditional.scala 39:67]
  wire  _GEN_250; // @[Conditional.scala 39:67]
  wire  _GEN_252; // @[Conditional.scala 39:67]
  wire  _GEN_253; // @[Conditional.scala 39:67]
  wire  _GEN_254; // @[Conditional.scala 39:67]
  wire  _GEN_255; // @[Conditional.scala 39:67]
  wire  _GEN_256; // @[Conditional.scala 39:67]
  wire  _GEN_257; // @[Conditional.scala 39:67]
  wire  _GEN_258; // @[Conditional.scala 39:67]
  wire  _GEN_259; // @[Conditional.scala 39:67]
  wire  _GEN_260; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_261; // @[Conditional.scala 39:67]
  wire  _GEN_262; // @[Conditional.scala 39:67]
  wire  _GEN_263; // @[Conditional.scala 39:67]
  wire  _GEN_265; // @[Conditional.scala 39:67]
  wire  _GEN_266; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_267; // @[Conditional.scala 39:67]
  wire  _GEN_268; // @[Conditional.scala 39:67]
  wire  _GEN_269; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_270; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_271; // @[Conditional.scala 39:67]
  wire  _GEN_272; // @[Conditional.scala 39:67]
  wire  _GEN_273; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_274; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_277; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_278; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_280; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_283; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_284; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_286; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_287; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_289; // @[Conditional.scala 39:67]
  wire  _GEN_292; // @[Conditional.scala 39:67]
  wire  _GEN_293; // @[Conditional.scala 39:67]
  wire  _GEN_294; // @[Conditional.scala 39:67]
  wire  _GEN_295; // @[Conditional.scala 39:67]
  wire  _GEN_296; // @[Conditional.scala 39:67]
  wire  _GEN_297; // @[Conditional.scala 39:67]
  wire  _GEN_298; // @[Conditional.scala 40:58]
  wire  _GEN_299; // @[Conditional.scala 40:58]
  wire  _GEN_300; // @[Conditional.scala 40:58]
  wire  _GEN_301; // @[Conditional.scala 40:58]
  wire  _GEN_302; // @[Conditional.scala 40:58]
  wire  _GEN_303; // @[Conditional.scala 40:58]
  wire  _GEN_304; // @[Conditional.scala 40:58]
  wire  _GEN_305; // @[Conditional.scala 40:58]
  wire  _GEN_306; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_307; // @[Conditional.scala 40:58]
  wire  _GEN_308; // @[Conditional.scala 40:58]
  wire  _GEN_309; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_310; // @[Conditional.scala 40:58]
  wire  _GEN_311; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_312; // @[Conditional.scala 40:58]
  wire  _GEN_313; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_314; // @[Conditional.scala 40:58]
  wire  _GEN_315; // @[Conditional.scala 40:58]
  wire  _GEN_316; // @[Conditional.scala 40:58]
  wire  _GEN_317; // @[Conditional.scala 40:58]
  wire  _GEN_318; // @[Conditional.scala 40:58]
  wire  _GEN_319; // @[Conditional.scala 40:58]
  wire  _GEN_320; // @[Conditional.scala 40:58]
  wire  _GEN_321; // @[Conditional.scala 40:58]
  wire  _GEN_322; // @[Conditional.scala 40:58]
  wire  _GEN_324; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_325; // @[Conditional.scala 40:58]
  wire  _GEN_326; // @[Conditional.scala 40:58]
  wire  _GEN_327; // @[Conditional.scala 40:58]
  wire  _GEN_329; // @[Conditional.scala 40:58]
  wire  _GEN_330; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_331; // @[Conditional.scala 40:58]
  wire  _GEN_332; // @[Conditional.scala 40:58]
  wire  _GEN_333; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_334; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_337; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_338; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_340; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_343; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_344; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_346; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_347; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_349; // @[Conditional.scala 40:58]
  wire  _GEN_352; // @[Conditional.scala 40:58]
  wire  _GEN_353; // @[Conditional.scala 40:58]
  wire  _GEN_354; // @[Conditional.scala 40:58]
  wire  _GEN_355; // @[Conditional.scala 40:58]
  wire  _GEN_356; // @[Conditional.scala 40:58]
  wire  _GEN_357; // @[Conditional.scala 40:58]
  assign _T_653 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_653 ? io_enable_bits_taskID : enable_R_taskID; // @[LoopBlock.scala 596:26]
  assign _GEN_2 = _T_653 ? io_enable_bits_control : enable_R_control; // @[LoopBlock.scala 596:26]
  assign _GEN_3 = _T_653 ? 1'h1 : enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_656 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_656 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_656 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_656 ? 1'h1 : loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_659 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_659 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_659 ? 1'h1 : loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_662 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_662 ? io_InLiveIn_0_bits_data : in_live_in_R_0_data; // @[LoopBlock.scala 623:33]
  assign _GEN_13 = _T_662 ? 1'h1 : in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_665 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_15 = _T_665 ? io_InLiveIn_1_bits_taskID : in_live_in_R_1_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_16 = _T_665 ? io_InLiveIn_1_bits_data : in_live_in_R_1_data; // @[LoopBlock.scala 623:33]
  assign _GEN_17 = _T_665 ? 1'h1 : in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_668 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_20 = _T_668 ? io_InLiveIn_2_bits_data : in_live_in_R_2_data; // @[LoopBlock.scala 623:33]
  assign _GEN_21 = _T_668 ? 1'h1 : in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_671 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_23 = _T_671 ? io_InLiveIn_3_bits_taskID : in_live_in_R_3_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_24 = _T_671 ? io_InLiveIn_3_bits_data : in_live_in_R_3_data; // @[LoopBlock.scala 623:33]
  assign _GEN_25 = _T_671 ? 1'h1 : in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_674 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_27 = _T_674 ? io_InLiveIn_4_bits_taskID : in_live_in_R_4_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_28 = _T_674 ? io_InLiveIn_4_bits_data : in_live_in_R_4_data; // @[LoopBlock.scala 623:33]
  assign _GEN_29 = _T_674 ? 1'h1 : in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_677 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 37:37]
  assign _GEN_32 = _T_677 ? io_InLiveIn_5_bits_data : in_live_in_R_5_data; // @[LoopBlock.scala 623:33]
  assign _GEN_33 = _T_677 ? 1'h1 : in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_680 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_35 = _T_680 ? io_CarryDepenIn_0_bits_taskID : in_carry_in_R_0_taskID; // @[LoopBlock.scala 641:37]
  assign _GEN_36 = _T_680 ? io_CarryDepenIn_0_bits_data : in_carry_in_R_0_data; // @[LoopBlock.scala 641:37]
  assign _GEN_37 = _T_680 ? 1'h1 : in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_682 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 37:37]
  assign _GEN_38 = _T_682 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_684 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 37:37]
  assign _GEN_39 = _T_684 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_686 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_40 = _T_686 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_41 = _T_686 ? 1'h1 : loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_689 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_42 = _T_689 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_43 = _T_689 ? 1'h1 : out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_692 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_44 = _T_692 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_45 = _T_692 ? 1'h1 : out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_695 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_46 = _T_695 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_47 = _T_695 ? 1'h1 : out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_698 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_48 = _T_698 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_49 = _T_698 ? 1'h1 : out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_701 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_50 = _T_701 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_51 = _T_701 ? 1'h1 : out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_704 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_52 = _T_704 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_53 = _T_704 ? 1'h1 : out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_707 = io_OutLiveIn_field5_1_ready & io_OutLiveIn_field5_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_54 = _T_707 ? 1'h0 : out_live_in_valid_R_5_1; // @[LoopBlock.scala 722:57]
  assign _GEN_55 = _T_707 ? 1'h1 : out_live_in_fire_R_5_1; // @[LoopBlock.scala 722:57]
  assign _T_710 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_56 = _T_710 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_714 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_715 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_716 = _T_715 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_717 = _T_716 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_718 = _T_717 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_719 = _T_718 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_720 = _T_719 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_58 = enable_R_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_59 = enable_R_control ? 1'h1 : _GEN_44; // @[LoopBlock.scala 870:26]
  assign _GEN_60 = enable_R_control ? 1'h1 : _GEN_46; // @[LoopBlock.scala 870:26]
  assign _GEN_61 = enable_R_control ? 1'h1 : _GEN_48; // @[LoopBlock.scala 870:26]
  assign _GEN_62 = enable_R_control ? 1'h1 : _GEN_50; // @[LoopBlock.scala 870:26]
  assign _GEN_63 = enable_R_control ? 1'h1 : _GEN_52; // @[LoopBlock.scala 870:26]
  assign _GEN_64 = enable_R_control ? 1'h1 : _GEN_54; // @[LoopBlock.scala 870:26]
  assign _GEN_65 = enable_R_control ? 1'h1 : _GEN_56; // @[LoopBlock.scala 870:26]
  assign _GEN_66 = enable_R_control ? 1'h1 : active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_67 = enable_R_control ? enable_R_taskID : active_loop_start_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_68 = enable_R_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_69 = enable_R_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_70 = enable_R_control ? enable_R_taskID : active_loop_back_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_71 = enable_R_control ? 1'h1 : _GEN_39; // @[LoopBlock.scala 870:26]
  assign _GEN_72 = enable_R_control ? 2'h1 : 2'h2; // @[LoopBlock.scala 870:26]
  assign _GEN_73 = enable_R_control ? loop_exit_R_0_control : 1'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_74 = enable_R_control ? loop_exit_R_0_taskID : 10'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_75 = enable_R_control ? _GEN_40 : 1'h1; // @[LoopBlock.scala 870:26]
  assign _GEN_76 = _T_720 ? _GEN_58 : _GEN_42; // @[LoopBlock.scala 869:48]
  assign _GEN_77 = _T_720 ? _GEN_59 : _GEN_44; // @[LoopBlock.scala 869:48]
  assign _GEN_78 = _T_720 ? _GEN_60 : _GEN_46; // @[LoopBlock.scala 869:48]
  assign _GEN_79 = _T_720 ? _GEN_61 : _GEN_48; // @[LoopBlock.scala 869:48]
  assign _GEN_80 = _T_720 ? _GEN_62 : _GEN_50; // @[LoopBlock.scala 869:48]
  assign _GEN_81 = _T_720 ? _GEN_63 : _GEN_52; // @[LoopBlock.scala 869:48]
  assign _GEN_82 = _T_720 ? _GEN_64 : _GEN_54; // @[LoopBlock.scala 869:48]
  assign _GEN_83 = _T_720 ? _GEN_65 : _GEN_56; // @[LoopBlock.scala 869:48]
  assign _GEN_84 = _T_720 ? _GEN_66 : active_loop_start_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_85 = _T_720 ? _GEN_67 : active_loop_start_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_86 = _T_720 ? _GEN_68 : _GEN_38; // @[LoopBlock.scala 869:48]
  assign _GEN_87 = _T_720 ? _GEN_69 : active_loop_back_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_88 = _T_720 ? _GEN_70 : active_loop_back_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_89 = _T_720 ? _GEN_71 : _GEN_39; // @[LoopBlock.scala 869:48]
  assign _GEN_90 = _T_720 ? _GEN_72 : state; // @[LoopBlock.scala 869:48]
  assign _GEN_91 = _T_720 ? _GEN_73 : loop_exit_R_0_control; // @[LoopBlock.scala 869:48]
  assign _GEN_92 = _T_720 ? _GEN_74 : loop_exit_R_0_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_93 = _T_720 ? _GEN_75 : _GEN_40; // @[LoopBlock.scala 869:48]
  assign _T_742 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_743 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_746 = out_live_in_fire_R_5_0 & out_live_in_fire_R_5_1; // @[LoopBlock.scala 825:65]
  assign _T_747 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_748 = _T_747 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_749 = _T_748 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_750 = _T_749 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_751 = _T_750 & _T_746; // @[LoopBlock.scala 828:26]
  assign _T_752 = _T_743 & _T_751; // @[LoopBlock.scala 899:29]
  assign _GEN_94 = loop_finish_R_0_control ? 1'h1 : _GEN_40; // @[LoopBlock.scala 936:64]
  assign _GEN_95 = loop_finish_R_0_control ? 1'h0 : active_loop_start_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_96 = loop_finish_R_0_control ? 10'h0 : active_loop_start_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_97 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_98 = loop_finish_R_0_control ? 10'h0 : active_loop_back_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_99 = loop_finish_R_0_control ? 1'h1 : loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_100 = loop_finish_R_0_control ? loop_back_R_0_taskID : loop_exit_R_0_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_101 = loop_finish_R_0_control ? 2'h2 : state; // @[LoopBlock.scala 936:64]
  assign _GEN_102 = loop_back_R_0_control ? 1'h0 : _GEN_95; // @[LoopBlock.scala 903:56]
  assign _GEN_103 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_96; // @[LoopBlock.scala 903:56]
  assign _GEN_104 = loop_back_R_0_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_105 = loop_back_R_0_control ? 1'h1 : _GEN_97; // @[LoopBlock.scala 903:56]
  assign _GEN_106 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_98; // @[LoopBlock.scala 903:56]
  assign _GEN_107 = loop_back_R_0_control ? 1'h1 : _GEN_39; // @[LoopBlock.scala 903:56]
  assign _GEN_108 = loop_back_R_0_control ? 1'h0 : _GEN_43; // @[LoopBlock.scala 903:56]
  assign _GEN_109 = loop_back_R_0_control ? 1'h0 : _GEN_45; // @[LoopBlock.scala 903:56]
  assign _GEN_110 = loop_back_R_0_control ? 1'h0 : _GEN_47; // @[LoopBlock.scala 903:56]
  assign _GEN_111 = loop_back_R_0_control ? 1'h0 : _GEN_49; // @[LoopBlock.scala 903:56]
  assign _GEN_112 = loop_back_R_0_control ? 1'h0 : _GEN_51; // @[LoopBlock.scala 903:56]
  assign _GEN_113 = loop_back_R_0_control ? 1'h0 : _GEN_53; // @[LoopBlock.scala 903:56]
  assign _GEN_114 = loop_back_R_0_control ? 1'h0 : _GEN_55; // @[LoopBlock.scala 903:56]
  assign _GEN_116 = loop_back_R_0_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_117 = loop_back_R_0_control ? 1'h1 : _GEN_44; // @[LoopBlock.scala 903:56]
  assign _GEN_118 = loop_back_R_0_control ? 1'h1 : _GEN_46; // @[LoopBlock.scala 903:56]
  assign _GEN_119 = loop_back_R_0_control ? 1'h1 : _GEN_48; // @[LoopBlock.scala 903:56]
  assign _GEN_120 = loop_back_R_0_control ? 1'h1 : _GEN_50; // @[LoopBlock.scala 903:56]
  assign _GEN_121 = loop_back_R_0_control ? 1'h1 : _GEN_52; // @[LoopBlock.scala 903:56]
  assign _GEN_122 = loop_back_R_0_control ? 1'h1 : _GEN_54; // @[LoopBlock.scala 903:56]
  assign _GEN_123 = loop_back_R_0_control ? 1'h1 : _GEN_56; // @[LoopBlock.scala 903:56]
  assign _GEN_124 = loop_back_R_0_control ? 1'h0 : _GEN_5; // @[LoopBlock.scala 903:56]
  assign _GEN_125 = loop_back_R_0_control ? 10'h0 : _GEN_4; // @[LoopBlock.scala 903:56]
  assign _GEN_126 = loop_back_R_0_control ? 1'h0 : _GEN_6; // @[LoopBlock.scala 903:56]
  assign _GEN_127 = loop_back_R_0_control ? 1'h0 : _GEN_8; // @[LoopBlock.scala 903:56]
  assign _GEN_129 = loop_back_R_0_control ? 1'h0 : _GEN_9; // @[LoopBlock.scala 903:56]
  assign _GEN_130 = loop_back_R_0_control ? 1'h0 : _GEN_37; // @[LoopBlock.scala 903:56]
  assign _GEN_131 = loop_back_R_0_control ? 2'h1 : _GEN_101; // @[LoopBlock.scala 903:56]
  assign _GEN_132 = loop_back_R_0_control ? _GEN_40 : _GEN_94; // @[LoopBlock.scala 903:56]
  assign _GEN_133 = loop_back_R_0_control ? loop_exit_R_0_control : _GEN_99; // @[LoopBlock.scala 903:56]
  assign _GEN_134 = loop_back_R_0_control ? loop_exit_R_0_taskID : _GEN_100; // @[LoopBlock.scala 903:56]
  assign _GEN_135 = _T_752 ? _GEN_102 : active_loop_start_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_136 = _T_752 ? _GEN_103 : active_loop_start_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_137 = _T_752 ? _GEN_104 : _GEN_38; // @[LoopBlock.scala 900:55]
  assign _GEN_138 = _T_752 ? _GEN_105 : active_loop_back_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_139 = _T_752 ? _GEN_106 : active_loop_back_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_140 = _T_752 ? _GEN_107 : _GEN_39; // @[LoopBlock.scala 900:55]
  assign _GEN_141 = _T_752 ? _GEN_108 : _GEN_43; // @[LoopBlock.scala 900:55]
  assign _GEN_142 = _T_752 ? _GEN_109 : _GEN_45; // @[LoopBlock.scala 900:55]
  assign _GEN_143 = _T_752 ? _GEN_110 : _GEN_47; // @[LoopBlock.scala 900:55]
  assign _GEN_144 = _T_752 ? _GEN_111 : _GEN_49; // @[LoopBlock.scala 900:55]
  assign _GEN_145 = _T_752 ? _GEN_112 : _GEN_51; // @[LoopBlock.scala 900:55]
  assign _GEN_146 = _T_752 ? _GEN_113 : _GEN_53; // @[LoopBlock.scala 900:55]
  assign _GEN_147 = _T_752 ? _GEN_114 : _GEN_55; // @[LoopBlock.scala 900:55]
  assign _GEN_149 = _T_752 ? _GEN_116 : _GEN_42; // @[LoopBlock.scala 900:55]
  assign _GEN_150 = _T_752 ? _GEN_117 : _GEN_44; // @[LoopBlock.scala 900:55]
  assign _GEN_151 = _T_752 ? _GEN_118 : _GEN_46; // @[LoopBlock.scala 900:55]
  assign _GEN_152 = _T_752 ? _GEN_119 : _GEN_48; // @[LoopBlock.scala 900:55]
  assign _GEN_153 = _T_752 ? _GEN_120 : _GEN_50; // @[LoopBlock.scala 900:55]
  assign _GEN_154 = _T_752 ? _GEN_121 : _GEN_52; // @[LoopBlock.scala 900:55]
  assign _GEN_155 = _T_752 ? _GEN_122 : _GEN_54; // @[LoopBlock.scala 900:55]
  assign _GEN_156 = _T_752 ? _GEN_123 : _GEN_56; // @[LoopBlock.scala 900:55]
  assign _GEN_157 = _T_752 ? _GEN_124 : _GEN_5; // @[LoopBlock.scala 900:55]
  assign _GEN_158 = _T_752 ? _GEN_125 : _GEN_4; // @[LoopBlock.scala 900:55]
  assign _GEN_159 = _T_752 ? _GEN_126 : _GEN_6; // @[LoopBlock.scala 900:55]
  assign _GEN_160 = _T_752 ? _GEN_127 : _GEN_8; // @[LoopBlock.scala 900:55]
  assign _GEN_162 = _T_752 ? _GEN_129 : _GEN_9; // @[LoopBlock.scala 900:55]
  assign _GEN_163 = _T_752 ? _GEN_130 : _GEN_37; // @[LoopBlock.scala 900:55]
  assign _GEN_164 = _T_752 ? _GEN_131 : state; // @[LoopBlock.scala 900:55]
  assign _GEN_165 = _T_752 ? _GEN_132 : _GEN_40; // @[LoopBlock.scala 900:55]
  assign _GEN_166 = _T_752 ? _GEN_133 : loop_exit_R_0_control; // @[LoopBlock.scala 900:55]
  assign _GEN_167 = _T_752 ? _GEN_134 : loop_exit_R_0_taskID; // @[LoopBlock.scala 900:55]
  assign _T_805 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_168 = loop_exit_fire_R_0 ? 10'h0 : _GEN_1; // @[LoopBlock.scala 955:48]
  assign _GEN_169 = loop_exit_fire_R_0 ? 1'h0 : _GEN_2; // @[LoopBlock.scala 955:48]
  assign _GEN_170 = loop_exit_fire_R_0 ? 1'h0 : _GEN_3; // @[LoopBlock.scala 955:48]
  assign _GEN_171 = loop_exit_fire_R_0 ? 1'h0 : _GEN_5; // @[LoopBlock.scala 955:48]
  assign _GEN_172 = loop_exit_fire_R_0 ? 10'h0 : _GEN_4; // @[LoopBlock.scala 955:48]
  assign _GEN_173 = loop_exit_fire_R_0 ? 1'h0 : _GEN_6; // @[LoopBlock.scala 955:48]
  assign _GEN_174 = loop_exit_fire_R_0 ? 1'h0 : _GEN_8; // @[LoopBlock.scala 955:48]
  assign _GEN_176 = loop_exit_fire_R_0 ? 1'h0 : _GEN_9; // @[LoopBlock.scala 955:48]
  assign _GEN_177 = loop_exit_fire_R_0 ? 32'h0 : _GEN_12; // @[LoopBlock.scala 955:48]
  assign _GEN_180 = loop_exit_fire_R_0 ? 32'h0 : _GEN_16; // @[LoopBlock.scala 955:48]
  assign _GEN_181 = loop_exit_fire_R_0 ? 10'h0 : _GEN_15; // @[LoopBlock.scala 955:48]
  assign _GEN_183 = loop_exit_fire_R_0 ? 32'h0 : _GEN_20; // @[LoopBlock.scala 955:48]
  assign _GEN_186 = loop_exit_fire_R_0 ? 32'h0 : _GEN_24; // @[LoopBlock.scala 955:48]
  assign _GEN_187 = loop_exit_fire_R_0 ? 10'h0 : _GEN_23; // @[LoopBlock.scala 955:48]
  assign _GEN_189 = loop_exit_fire_R_0 ? 32'h0 : _GEN_28; // @[LoopBlock.scala 955:48]
  assign _GEN_190 = loop_exit_fire_R_0 ? 10'h0 : _GEN_27; // @[LoopBlock.scala 955:48]
  assign _GEN_192 = loop_exit_fire_R_0 ? 32'h0 : _GEN_32; // @[LoopBlock.scala 955:48]
  assign _GEN_195 = loop_exit_fire_R_0 ? 1'h0 : _GEN_13; // @[LoopBlock.scala 955:48]
  assign _GEN_196 = loop_exit_fire_R_0 ? 1'h0 : _GEN_17; // @[LoopBlock.scala 955:48]
  assign _GEN_197 = loop_exit_fire_R_0 ? 1'h0 : _GEN_21; // @[LoopBlock.scala 955:48]
  assign _GEN_198 = loop_exit_fire_R_0 ? 1'h0 : _GEN_25; // @[LoopBlock.scala 955:48]
  assign _GEN_199 = loop_exit_fire_R_0 ? 1'h0 : _GEN_29; // @[LoopBlock.scala 955:48]
  assign _GEN_200 = loop_exit_fire_R_0 ? 1'h0 : _GEN_33; // @[LoopBlock.scala 955:48]
  assign _GEN_201 = loop_exit_fire_R_0 ? 1'h0 : _GEN_37; // @[LoopBlock.scala 955:48]
  assign _GEN_202 = loop_exit_fire_R_0 ? 2'h0 : state; // @[LoopBlock.scala 955:48]
  assign _GEN_203 = _T_805 ? _GEN_168 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_204 = _T_805 ? _GEN_169 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_205 = _T_805 ? _GEN_170 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_206 = _T_805 ? _GEN_171 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_207 = _T_805 ? _GEN_172 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_208 = _T_805 ? _GEN_173 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_209 = _T_805 ? _GEN_174 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_211 = _T_805 ? _GEN_176 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_212 = _T_805 ? _GEN_177 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_215 = _T_805 ? _GEN_180 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_216 = _T_805 ? _GEN_181 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_218 = _T_805 ? _GEN_183 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_221 = _T_805 ? _GEN_186 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_222 = _T_805 ? _GEN_187 : _GEN_23; // @[Conditional.scala 39:67]
  assign _GEN_224 = _T_805 ? _GEN_189 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_225 = _T_805 ? _GEN_190 : _GEN_27; // @[Conditional.scala 39:67]
  assign _GEN_227 = _T_805 ? _GEN_192 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_230 = _T_805 ? _GEN_195 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_231 = _T_805 ? _GEN_196 : _GEN_17; // @[Conditional.scala 39:67]
  assign _GEN_232 = _T_805 ? _GEN_197 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_233 = _T_805 ? _GEN_198 : _GEN_25; // @[Conditional.scala 39:67]
  assign _GEN_234 = _T_805 ? _GEN_199 : _GEN_29; // @[Conditional.scala 39:67]
  assign _GEN_235 = _T_805 ? _GEN_200 : _GEN_33; // @[Conditional.scala 39:67]
  assign _GEN_236 = _T_805 ? _GEN_201 : _GEN_37; // @[Conditional.scala 39:67]
  assign _GEN_237 = _T_805 ? _GEN_202 : state; // @[Conditional.scala 39:67]
  assign _GEN_238 = _T_742 ? _GEN_135 : active_loop_start_R_control; // @[Conditional.scala 39:67]
  assign _GEN_239 = _T_742 ? _GEN_136 : active_loop_start_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_240 = _T_742 ? _GEN_137 : _GEN_38; // @[Conditional.scala 39:67]
  assign _GEN_241 = _T_742 ? _GEN_138 : active_loop_back_R_control; // @[Conditional.scala 39:67]
  assign _GEN_242 = _T_742 ? _GEN_139 : active_loop_back_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_243 = _T_742 ? _GEN_140 : _GEN_39; // @[Conditional.scala 39:67]
  assign _GEN_244 = _T_742 ? _GEN_141 : _GEN_43; // @[Conditional.scala 39:67]
  assign _GEN_245 = _T_742 ? _GEN_142 : _GEN_45; // @[Conditional.scala 39:67]
  assign _GEN_246 = _T_742 ? _GEN_143 : _GEN_47; // @[Conditional.scala 39:67]
  assign _GEN_247 = _T_742 ? _GEN_144 : _GEN_49; // @[Conditional.scala 39:67]
  assign _GEN_248 = _T_742 ? _GEN_145 : _GEN_51; // @[Conditional.scala 39:67]
  assign _GEN_249 = _T_742 ? _GEN_146 : _GEN_53; // @[Conditional.scala 39:67]
  assign _GEN_250 = _T_742 ? _GEN_147 : _GEN_55; // @[Conditional.scala 39:67]
  assign _GEN_252 = _T_742 ? _GEN_149 : _GEN_42; // @[Conditional.scala 39:67]
  assign _GEN_253 = _T_742 ? _GEN_150 : _GEN_44; // @[Conditional.scala 39:67]
  assign _GEN_254 = _T_742 ? _GEN_151 : _GEN_46; // @[Conditional.scala 39:67]
  assign _GEN_255 = _T_742 ? _GEN_152 : _GEN_48; // @[Conditional.scala 39:67]
  assign _GEN_256 = _T_742 ? _GEN_153 : _GEN_50; // @[Conditional.scala 39:67]
  assign _GEN_257 = _T_742 ? _GEN_154 : _GEN_52; // @[Conditional.scala 39:67]
  assign _GEN_258 = _T_742 ? _GEN_155 : _GEN_54; // @[Conditional.scala 39:67]
  assign _GEN_259 = _T_742 ? _GEN_156 : _GEN_56; // @[Conditional.scala 39:67]
  assign _GEN_260 = _T_742 ? _GEN_157 : _GEN_206; // @[Conditional.scala 39:67]
  assign _GEN_261 = _T_742 ? _GEN_158 : _GEN_207; // @[Conditional.scala 39:67]
  assign _GEN_262 = _T_742 ? _GEN_159 : _GEN_208; // @[Conditional.scala 39:67]
  assign _GEN_263 = _T_742 ? _GEN_160 : _GEN_209; // @[Conditional.scala 39:67]
  assign _GEN_265 = _T_742 ? _GEN_162 : _GEN_211; // @[Conditional.scala 39:67]
  assign _GEN_266 = _T_742 ? _GEN_163 : _GEN_236; // @[Conditional.scala 39:67]
  assign _GEN_267 = _T_742 ? _GEN_164 : _GEN_237; // @[Conditional.scala 39:67]
  assign _GEN_268 = _T_742 ? _GEN_165 : _GEN_40; // @[Conditional.scala 39:67]
  assign _GEN_269 = _T_742 ? _GEN_166 : loop_exit_R_0_control; // @[Conditional.scala 39:67]
  assign _GEN_270 = _T_742 ? _GEN_167 : loop_exit_R_0_taskID; // @[Conditional.scala 39:67]
  assign _GEN_271 = _T_742 ? _GEN_1 : _GEN_203; // @[Conditional.scala 39:67]
  assign _GEN_272 = _T_742 ? _GEN_2 : _GEN_204; // @[Conditional.scala 39:67]
  assign _GEN_273 = _T_742 ? _GEN_3 : _GEN_205; // @[Conditional.scala 39:67]
  assign _GEN_274 = _T_742 ? _GEN_12 : _GEN_212; // @[Conditional.scala 39:67]
  assign _GEN_277 = _T_742 ? _GEN_16 : _GEN_215; // @[Conditional.scala 39:67]
  assign _GEN_278 = _T_742 ? _GEN_15 : _GEN_216; // @[Conditional.scala 39:67]
  assign _GEN_280 = _T_742 ? _GEN_20 : _GEN_218; // @[Conditional.scala 39:67]
  assign _GEN_283 = _T_742 ? _GEN_24 : _GEN_221; // @[Conditional.scala 39:67]
  assign _GEN_284 = _T_742 ? _GEN_23 : _GEN_222; // @[Conditional.scala 39:67]
  assign _GEN_286 = _T_742 ? _GEN_28 : _GEN_224; // @[Conditional.scala 39:67]
  assign _GEN_287 = _T_742 ? _GEN_27 : _GEN_225; // @[Conditional.scala 39:67]
  assign _GEN_289 = _T_742 ? _GEN_32 : _GEN_227; // @[Conditional.scala 39:67]
  assign _GEN_292 = _T_742 ? _GEN_13 : _GEN_230; // @[Conditional.scala 39:67]
  assign _GEN_293 = _T_742 ? _GEN_17 : _GEN_231; // @[Conditional.scala 39:67]
  assign _GEN_294 = _T_742 ? _GEN_21 : _GEN_232; // @[Conditional.scala 39:67]
  assign _GEN_295 = _T_742 ? _GEN_25 : _GEN_233; // @[Conditional.scala 39:67]
  assign _GEN_296 = _T_742 ? _GEN_29 : _GEN_234; // @[Conditional.scala 39:67]
  assign _GEN_297 = _T_742 ? _GEN_33 : _GEN_235; // @[Conditional.scala 39:67]
  assign _GEN_298 = _T_714 ? _GEN_76 : _GEN_252; // @[Conditional.scala 40:58]
  assign _GEN_299 = _T_714 ? _GEN_77 : _GEN_253; // @[Conditional.scala 40:58]
  assign _GEN_300 = _T_714 ? _GEN_78 : _GEN_254; // @[Conditional.scala 40:58]
  assign _GEN_301 = _T_714 ? _GEN_79 : _GEN_255; // @[Conditional.scala 40:58]
  assign _GEN_302 = _T_714 ? _GEN_80 : _GEN_256; // @[Conditional.scala 40:58]
  assign _GEN_303 = _T_714 ? _GEN_81 : _GEN_257; // @[Conditional.scala 40:58]
  assign _GEN_304 = _T_714 ? _GEN_82 : _GEN_258; // @[Conditional.scala 40:58]
  assign _GEN_305 = _T_714 ? _GEN_83 : _GEN_259; // @[Conditional.scala 40:58]
  assign _GEN_306 = _T_714 ? _GEN_84 : _GEN_238; // @[Conditional.scala 40:58]
  assign _GEN_307 = _T_714 ? _GEN_85 : _GEN_239; // @[Conditional.scala 40:58]
  assign _GEN_308 = _T_714 ? _GEN_86 : _GEN_240; // @[Conditional.scala 40:58]
  assign _GEN_309 = _T_714 ? _GEN_87 : _GEN_241; // @[Conditional.scala 40:58]
  assign _GEN_310 = _T_714 ? _GEN_88 : _GEN_242; // @[Conditional.scala 40:58]
  assign _GEN_311 = _T_714 ? _GEN_89 : _GEN_243; // @[Conditional.scala 40:58]
  assign _GEN_312 = _T_714 ? _GEN_90 : _GEN_267; // @[Conditional.scala 40:58]
  assign _GEN_313 = _T_714 ? _GEN_91 : _GEN_269; // @[Conditional.scala 40:58]
  assign _GEN_314 = _T_714 ? _GEN_92 : _GEN_270; // @[Conditional.scala 40:58]
  assign _GEN_315 = _T_714 ? _GEN_93 : _GEN_268; // @[Conditional.scala 40:58]
  assign _GEN_316 = _T_714 ? _GEN_43 : _GEN_244; // @[Conditional.scala 40:58]
  assign _GEN_317 = _T_714 ? _GEN_45 : _GEN_245; // @[Conditional.scala 40:58]
  assign _GEN_318 = _T_714 ? _GEN_47 : _GEN_246; // @[Conditional.scala 40:58]
  assign _GEN_319 = _T_714 ? _GEN_49 : _GEN_247; // @[Conditional.scala 40:58]
  assign _GEN_320 = _T_714 ? _GEN_51 : _GEN_248; // @[Conditional.scala 40:58]
  assign _GEN_321 = _T_714 ? _GEN_53 : _GEN_249; // @[Conditional.scala 40:58]
  assign _GEN_322 = _T_714 ? _GEN_55 : _GEN_250; // @[Conditional.scala 40:58]
  assign _GEN_324 = _T_714 ? _GEN_5 : _GEN_260; // @[Conditional.scala 40:58]
  assign _GEN_325 = _T_714 ? _GEN_4 : _GEN_261; // @[Conditional.scala 40:58]
  assign _GEN_326 = _T_714 ? _GEN_6 : _GEN_262; // @[Conditional.scala 40:58]
  assign _GEN_327 = _T_714 ? _GEN_8 : _GEN_263; // @[Conditional.scala 40:58]
  assign _GEN_329 = _T_714 ? _GEN_9 : _GEN_265; // @[Conditional.scala 40:58]
  assign _GEN_330 = _T_714 ? _GEN_37 : _GEN_266; // @[Conditional.scala 40:58]
  assign _GEN_331 = _T_714 ? _GEN_1 : _GEN_271; // @[Conditional.scala 40:58]
  assign _GEN_332 = _T_714 ? _GEN_2 : _GEN_272; // @[Conditional.scala 40:58]
  assign _GEN_333 = _T_714 ? _GEN_3 : _GEN_273; // @[Conditional.scala 40:58]
  assign _GEN_334 = _T_714 ? _GEN_12 : _GEN_274; // @[Conditional.scala 40:58]
  assign _GEN_337 = _T_714 ? _GEN_16 : _GEN_277; // @[Conditional.scala 40:58]
  assign _GEN_338 = _T_714 ? _GEN_15 : _GEN_278; // @[Conditional.scala 40:58]
  assign _GEN_340 = _T_714 ? _GEN_20 : _GEN_280; // @[Conditional.scala 40:58]
  assign _GEN_343 = _T_714 ? _GEN_24 : _GEN_283; // @[Conditional.scala 40:58]
  assign _GEN_344 = _T_714 ? _GEN_23 : _GEN_284; // @[Conditional.scala 40:58]
  assign _GEN_346 = _T_714 ? _GEN_28 : _GEN_286; // @[Conditional.scala 40:58]
  assign _GEN_347 = _T_714 ? _GEN_27 : _GEN_287; // @[Conditional.scala 40:58]
  assign _GEN_349 = _T_714 ? _GEN_32 : _GEN_289; // @[Conditional.scala 40:58]
  assign _GEN_352 = _T_714 ? _GEN_13 : _GEN_292; // @[Conditional.scala 40:58]
  assign _GEN_353 = _T_714 ? _GEN_17 : _GEN_293; // @[Conditional.scala 40:58]
  assign _GEN_354 = _T_714 ? _GEN_21 : _GEN_294; // @[Conditional.scala 40:58]
  assign _GEN_355 = _T_714 ? _GEN_25 : _GEN_295; // @[Conditional.scala 40:58]
  assign _GEN_356 = _T_714 ? _GEN_29 : _GEN_296; // @[Conditional.scala 40:58]
  assign _GEN_357 = _T_714 ? _GEN_33 : _GEN_297; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_1_valid = out_live_in_valid_R_5_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_1_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_taskID = in_live_in_R_3_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_3_taskID = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_14[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_23[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_live_in_valid_R_5_1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  out_live_in_fire_R_5_1 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_41[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_44[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_47[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  state = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_653) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_742) begin
          if (_T_653) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_653) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_653) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_653) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_742) begin
          if (_T_653) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_653) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_653) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_653) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_653) begin
            enable_valid_R <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_653) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_653) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_656) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_656) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_656) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_656) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_656) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_656) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_656) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_656) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_656) begin
          loop_back_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_656) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_656) begin
              loop_back_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_656) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_659) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_659) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_659) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_659) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_8;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_659) begin
          loop_finish_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_659) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_659) begin
              loop_finish_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_659) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_714) begin
        if (_T_662) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_742) begin
          if (_T_662) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_662) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_662) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_665) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_742) begin
          if (_T_665) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_taskID <= 10'h0;
            end else begin
              if (_T_665) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_665) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_714) begin
        if (_T_665) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_742) begin
          if (_T_665) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_665) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_665) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_714) begin
        if (_T_668) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_742) begin
          if (_T_668) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_668) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_668) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_671) begin
          in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
        end
      end else begin
        if (_T_742) begin
          if (_T_671) begin
            in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_taskID <= 10'h0;
            end else begin
              if (_T_671) begin
                in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
              end
            end
          end else begin
            if (_T_671) begin
              in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_714) begin
        if (_T_671) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_742) begin
          if (_T_671) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_671) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_671) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_674) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_742) begin
          if (_T_674) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 10'h0;
            end else begin
              if (_T_674) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_674) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_714) begin
        if (_T_674) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_742) begin
          if (_T_674) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_674) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_674) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_714) begin
        if (_T_677) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_742) begin
          if (_T_677) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_677) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_677) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_662) begin
          in_live_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_662) begin
            in_live_in_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_662) begin
                in_live_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_662) begin
              in_live_in_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_665) begin
          in_live_in_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_665) begin
            in_live_in_valid_R_1 <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              if (_T_665) begin
                in_live_in_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_665) begin
              in_live_in_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_668) begin
          in_live_in_valid_R_2 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_668) begin
            in_live_in_valid_R_2 <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              if (_T_668) begin
                in_live_in_valid_R_2 <= 1'h1;
              end
            end
          end else begin
            if (_T_668) begin
              in_live_in_valid_R_2 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_671) begin
          in_live_in_valid_R_3 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_671) begin
            in_live_in_valid_R_3 <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              if (_T_671) begin
                in_live_in_valid_R_3 <= 1'h1;
              end
            end
          end else begin
            if (_T_671) begin
              in_live_in_valid_R_3 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_674) begin
          in_live_in_valid_R_4 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_674) begin
            in_live_in_valid_R_4 <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              if (_T_674) begin
                in_live_in_valid_R_4 <= 1'h1;
              end
            end
          end else begin
            if (_T_674) begin
              in_live_in_valid_R_4 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_677) begin
          in_live_in_valid_R_5 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_677) begin
            in_live_in_valid_R_5 <= 1'h1;
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              if (_T_677) begin
                in_live_in_valid_R_5 <= 1'h1;
              end
            end
          end else begin
            if (_T_677) begin
              in_live_in_valid_R_5 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_680) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_680) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_680) begin
          in_carry_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_680) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_680) begin
              in_carry_in_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_680) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_689) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_689) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_689) begin
                out_live_in_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_689) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_0_0 <= _GEN_42;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_1_0 <= 1'h1;
          end else begin
            if (_T_692) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_692) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_1_0 <= 1'h1;
            end else begin
              if (_T_692) begin
                out_live_in_valid_R_1_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_692) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_1_0 <= _GEN_44;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_2_0 <= 1'h1;
          end else begin
            if (_T_695) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_695) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_2_0 <= 1'h1;
            end else begin
              if (_T_695) begin
                out_live_in_valid_R_2_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_695) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_2_0 <= _GEN_46;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_3_0 <= 1'h1;
          end else begin
            if (_T_698) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_698) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_3_0 <= 1'h1;
            end else begin
              if (_T_698) begin
                out_live_in_valid_R_3_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_698) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_3_0 <= _GEN_48;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_4_0 <= 1'h1;
          end else begin
            if (_T_701) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_701) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_4_0 <= 1'h1;
            end else begin
              if (_T_701) begin
                out_live_in_valid_R_4_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_701) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_4_0 <= _GEN_50;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_5_0 <= 1'h1;
          end else begin
            if (_T_704) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_704) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_5_0 <= 1'h1;
            end else begin
              if (_T_704) begin
                out_live_in_valid_R_5_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_704) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_5_0 <= _GEN_52;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_1 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_live_in_valid_R_5_1 <= 1'h1;
          end else begin
            if (_T_707) begin
              out_live_in_valid_R_5_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_707) begin
            out_live_in_valid_R_5_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_5_1 <= 1'h1;
            end else begin
              if (_T_707) begin
                out_live_in_valid_R_5_1 <= 1'h0;
              end
            end
          end else begin
            if (_T_707) begin
              out_live_in_valid_R_5_1 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_5_1 <= _GEN_54;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_689) begin
          out_live_in_fire_R_0_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              if (_T_689) begin
                out_live_in_fire_R_0_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_689) begin
              out_live_in_fire_R_0_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_689) begin
            out_live_in_fire_R_0_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_692) begin
          out_live_in_fire_R_1_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              if (_T_692) begin
                out_live_in_fire_R_1_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_692) begin
              out_live_in_fire_R_1_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_692) begin
            out_live_in_fire_R_1_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_695) begin
          out_live_in_fire_R_2_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              if (_T_695) begin
                out_live_in_fire_R_2_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_695) begin
              out_live_in_fire_R_2_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_695) begin
            out_live_in_fire_R_2_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_698) begin
          out_live_in_fire_R_3_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              if (_T_698) begin
                out_live_in_fire_R_3_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_698) begin
              out_live_in_fire_R_3_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_698) begin
            out_live_in_fire_R_3_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_701) begin
          out_live_in_fire_R_4_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              if (_T_701) begin
                out_live_in_fire_R_4_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_701) begin
              out_live_in_fire_R_4_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_701) begin
            out_live_in_fire_R_4_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_704) begin
          out_live_in_fire_R_5_0 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              if (_T_704) begin
                out_live_in_fire_R_5_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_704) begin
              out_live_in_fire_R_5_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_704) begin
            out_live_in_fire_R_5_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_1 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_707) begin
          out_live_in_fire_R_5_1 <= 1'h1;
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_1 <= 1'h0;
            end else begin
              if (_T_707) begin
                out_live_in_fire_R_5_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_707) begin
              out_live_in_fire_R_5_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_707) begin
            out_live_in_fire_R_5_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            out_carry_out_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_710) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_710) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              out_carry_out_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_710) begin
                out_carry_out_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_710) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_carry_out_valid_R_0_0 <= _GEN_56;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            active_loop_start_R_control <= 1'h1;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            active_loop_start_valid_R <= 1'h1;
          end else begin
            if (_T_682) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_682) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              active_loop_start_valid_R <= 1'h1;
            end else begin
              if (_T_682) begin
                active_loop_start_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_682) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_start_valid_R <= _GEN_38;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_control <= 1'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            active_loop_back_valid_R <= 1'h1;
          end else begin
            if (_T_684) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_684) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              active_loop_back_valid_R <= 1'h1;
            end else begin
              if (_T_684) begin
                active_loop_back_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_684) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_back_valid_R <= _GEN_39;
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 10'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 10'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_control <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_control <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            if (_T_686) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_686) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              if (_T_686) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              if (loop_finish_R_0_control) begin
                loop_exit_valid_R_0 <= 1'h1;
              end else begin
                if (_T_686) begin
                  loop_exit_valid_R_0 <= 1'h0;
                end
              end
            end
          end else begin
            loop_exit_valid_R_0 <= _GEN_40;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      if (_T_686) begin
        loop_exit_fire_R_0 <= 1'h1;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_714) begin
        if (_T_720) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_742) begin
          if (_T_752) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_805) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [9:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [9:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [9:0]  io_InLiveIn_5_bits_taskID,
  input  [31:0] io_InLiveIn_5_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [9:0]  io_OutLiveIn_field5_0_bits_taskID,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field4_1_ready,
  output        io_OutLiveIn_field4_1_valid,
  output [31:0] io_OutLiveIn_field4_1_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [9:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [9:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_OutLiveIn_field0_1_ready,
  output        io_OutLiveIn_field0_1_valid,
  output [31:0] io_OutLiveIn_field0_1_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [9:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [9:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [9:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [9:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [9:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [9:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_2;
  reg [9:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_3;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_5;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_6;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_7;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_8;
  reg [9:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [9:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [9:0] in_live_in_R_5_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_17;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_18;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_19;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_20;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_21;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_22;
  reg [9:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_23;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_24;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_25;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_26;
  reg  out_live_in_valid_R_0_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_29;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_30;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_31;
  reg  out_live_in_valid_R_4_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_32;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_33;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_34;
  reg  out_live_in_fire_R_0_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_35;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_36;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_37;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_38;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_39;
  reg  out_live_in_fire_R_4_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_40;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_41;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_42;
  reg [9:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_43;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_44;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_45;
  reg [9:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_46;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_47;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_48;
  reg [9:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_49;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_50;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_51;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_52;
  wire  _T_671; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[LoopBlock.scala 596:26]
  wire  _GEN_2; // @[LoopBlock.scala 596:26]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_674; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_4; // @[LoopBlock.scala 603:33]
  wire  _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_677; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_680; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[LoopBlock.scala 623:33]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_683; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_15; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_16; // @[LoopBlock.scala 623:33]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_686; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_19; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_20; // @[LoopBlock.scala 623:33]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_689; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_24; // @[LoopBlock.scala 623:33]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_692; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_28; // @[LoopBlock.scala 623:33]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_695; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_31; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_32; // @[LoopBlock.scala 623:33]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_698; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_35; // @[LoopBlock.scala 641:37]
  wire [31:0] _GEN_36; // @[LoopBlock.scala 641:37]
  wire  _GEN_37; // @[LoopBlock.scala 641:37]
  wire  _T_700; // @[Decoupled.scala 37:37]
  wire  _GEN_38; // @[LoopBlock.scala 704:39]
  wire  _T_702; // @[Decoupled.scala 37:37]
  wire  _GEN_39; // @[LoopBlock.scala 708:38]
  wire  _T_704; // @[Decoupled.scala 37:37]
  wire  _GEN_40; // @[LoopBlock.scala 713:33]
  wire  _GEN_41; // @[LoopBlock.scala 713:33]
  wire  _T_707; // @[Decoupled.scala 37:37]
  wire  _GEN_42; // @[LoopBlock.scala 722:57]
  wire  _GEN_43; // @[LoopBlock.scala 722:57]
  wire  _T_710; // @[Decoupled.scala 37:37]
  wire  _GEN_44; // @[LoopBlock.scala 722:57]
  wire  _GEN_45; // @[LoopBlock.scala 722:57]
  wire  _T_713; // @[Decoupled.scala 37:37]
  wire  _GEN_46; // @[LoopBlock.scala 722:57]
  wire  _GEN_47; // @[LoopBlock.scala 722:57]
  wire  _T_716; // @[Decoupled.scala 37:37]
  wire  _GEN_48; // @[LoopBlock.scala 722:57]
  wire  _GEN_49; // @[LoopBlock.scala 722:57]
  wire  _T_719; // @[Decoupled.scala 37:37]
  wire  _GEN_50; // @[LoopBlock.scala 722:57]
  wire  _GEN_51; // @[LoopBlock.scala 722:57]
  wire  _T_722; // @[Decoupled.scala 37:37]
  wire  _GEN_52; // @[LoopBlock.scala 722:57]
  wire  _GEN_53; // @[LoopBlock.scala 722:57]
  wire  _T_725; // @[Decoupled.scala 37:37]
  wire  _GEN_54; // @[LoopBlock.scala 722:57]
  wire  _GEN_55; // @[LoopBlock.scala 722:57]
  wire  _T_728; // @[Decoupled.scala 37:37]
  wire  _GEN_56; // @[LoopBlock.scala 722:57]
  wire  _GEN_57; // @[LoopBlock.scala 722:57]
  wire  _T_731; // @[Decoupled.scala 37:37]
  wire  _GEN_58; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_53;
  wire  _T_735; // @[Conditional.scala 37:30]
  wire  _T_736; // @[LoopBlock.scala 765:35]
  wire  _T_737; // @[LoopBlock.scala 765:35]
  wire  _T_738; // @[LoopBlock.scala 765:35]
  wire  _T_739; // @[LoopBlock.scala 765:35]
  wire  _T_740; // @[LoopBlock.scala 765:35]
  wire  _T_741; // @[LoopBlock.scala 869:28]
  wire  _GEN_60; // @[LoopBlock.scala 870:26]
  wire  _GEN_61; // @[LoopBlock.scala 870:26]
  wire  _GEN_62; // @[LoopBlock.scala 870:26]
  wire  _GEN_63; // @[LoopBlock.scala 870:26]
  wire  _GEN_64; // @[LoopBlock.scala 870:26]
  wire  _GEN_65; // @[LoopBlock.scala 870:26]
  wire  _GEN_66; // @[LoopBlock.scala 870:26]
  wire  _GEN_67; // @[LoopBlock.scala 870:26]
  wire  _GEN_68; // @[LoopBlock.scala 870:26]
  wire  _GEN_69; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_70; // @[LoopBlock.scala 870:26]
  wire  _GEN_71; // @[LoopBlock.scala 870:26]
  wire  _GEN_72; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_73; // @[LoopBlock.scala 870:26]
  wire  _GEN_74; // @[LoopBlock.scala 870:26]
  wire [1:0] _GEN_75; // @[LoopBlock.scala 870:26]
  wire  _GEN_76; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_77; // @[LoopBlock.scala 870:26]
  wire  _GEN_78; // @[LoopBlock.scala 870:26]
  wire  _GEN_79; // @[LoopBlock.scala 869:48]
  wire  _GEN_80; // @[LoopBlock.scala 869:48]
  wire  _GEN_81; // @[LoopBlock.scala 869:48]
  wire  _GEN_82; // @[LoopBlock.scala 869:48]
  wire  _GEN_83; // @[LoopBlock.scala 869:48]
  wire  _GEN_84; // @[LoopBlock.scala 869:48]
  wire  _GEN_85; // @[LoopBlock.scala 869:48]
  wire  _GEN_86; // @[LoopBlock.scala 869:48]
  wire  _GEN_87; // @[LoopBlock.scala 869:48]
  wire  _GEN_88; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_89; // @[LoopBlock.scala 869:48]
  wire  _GEN_90; // @[LoopBlock.scala 869:48]
  wire  _GEN_91; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_92; // @[LoopBlock.scala 869:48]
  wire  _GEN_93; // @[LoopBlock.scala 869:48]
  wire [1:0] _GEN_94; // @[LoopBlock.scala 869:48]
  wire  _GEN_95; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_96; // @[LoopBlock.scala 869:48]
  wire  _GEN_97; // @[LoopBlock.scala 869:48]
  wire  _T_764; // @[Conditional.scala 37:30]
  wire  _T_765; // @[LoopBlock.scala 898:30]
  wire  _T_768; // @[LoopBlock.scala 825:65]
  wire  _T_769; // @[LoopBlock.scala 825:65]
  wire  _T_770; // @[LoopBlock.scala 828:26]
  wire  _T_771; // @[LoopBlock.scala 828:26]
  wire  _T_772; // @[LoopBlock.scala 828:26]
  wire  _T_773; // @[LoopBlock.scala 828:26]
  wire  _T_774; // @[LoopBlock.scala 828:26]
  wire  _T_775; // @[LoopBlock.scala 899:29]
  wire  _GEN_98; // @[LoopBlock.scala 936:64]
  wire  _GEN_99; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_100; // @[LoopBlock.scala 936:64]
  wire  _GEN_101; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_102; // @[LoopBlock.scala 936:64]
  wire  _GEN_103; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_104; // @[LoopBlock.scala 936:64]
  wire [1:0] _GEN_105; // @[LoopBlock.scala 936:64]
  wire  _GEN_106; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_107; // @[LoopBlock.scala 903:56]
  wire  _GEN_108; // @[LoopBlock.scala 903:56]
  wire  _GEN_109; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_110; // @[LoopBlock.scala 903:56]
  wire  _GEN_111; // @[LoopBlock.scala 903:56]
  wire  _GEN_112; // @[LoopBlock.scala 903:56]
  wire  _GEN_113; // @[LoopBlock.scala 903:56]
  wire  _GEN_114; // @[LoopBlock.scala 903:56]
  wire  _GEN_115; // @[LoopBlock.scala 903:56]
  wire  _GEN_116; // @[LoopBlock.scala 903:56]
  wire  _GEN_117; // @[LoopBlock.scala 903:56]
  wire  _GEN_118; // @[LoopBlock.scala 903:56]
  wire  _GEN_119; // @[LoopBlock.scala 903:56]
  wire  _GEN_121; // @[LoopBlock.scala 903:56]
  wire  _GEN_122; // @[LoopBlock.scala 903:56]
  wire  _GEN_123; // @[LoopBlock.scala 903:56]
  wire  _GEN_124; // @[LoopBlock.scala 903:56]
  wire  _GEN_125; // @[LoopBlock.scala 903:56]
  wire  _GEN_126; // @[LoopBlock.scala 903:56]
  wire  _GEN_127; // @[LoopBlock.scala 903:56]
  wire  _GEN_128; // @[LoopBlock.scala 903:56]
  wire  _GEN_129; // @[LoopBlock.scala 903:56]
  wire  _GEN_130; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_131; // @[LoopBlock.scala 903:56]
  wire  _GEN_132; // @[LoopBlock.scala 903:56]
  wire  _GEN_133; // @[LoopBlock.scala 903:56]
  wire  _GEN_135; // @[LoopBlock.scala 903:56]
  wire  _GEN_136; // @[LoopBlock.scala 903:56]
  wire [1:0] _GEN_137; // @[LoopBlock.scala 903:56]
  wire  _GEN_138; // @[LoopBlock.scala 903:56]
  wire  _GEN_139; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_140; // @[LoopBlock.scala 903:56]
  wire  _GEN_141; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_142; // @[LoopBlock.scala 900:55]
  wire  _GEN_143; // @[LoopBlock.scala 900:55]
  wire  _GEN_144; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_145; // @[LoopBlock.scala 900:55]
  wire  _GEN_146; // @[LoopBlock.scala 900:55]
  wire  _GEN_147; // @[LoopBlock.scala 900:55]
  wire  _GEN_148; // @[LoopBlock.scala 900:55]
  wire  _GEN_149; // @[LoopBlock.scala 900:55]
  wire  _GEN_150; // @[LoopBlock.scala 900:55]
  wire  _GEN_151; // @[LoopBlock.scala 900:55]
  wire  _GEN_152; // @[LoopBlock.scala 900:55]
  wire  _GEN_153; // @[LoopBlock.scala 900:55]
  wire  _GEN_154; // @[LoopBlock.scala 900:55]
  wire  _GEN_156; // @[LoopBlock.scala 900:55]
  wire  _GEN_157; // @[LoopBlock.scala 900:55]
  wire  _GEN_158; // @[LoopBlock.scala 900:55]
  wire  _GEN_159; // @[LoopBlock.scala 900:55]
  wire  _GEN_160; // @[LoopBlock.scala 900:55]
  wire  _GEN_161; // @[LoopBlock.scala 900:55]
  wire  _GEN_162; // @[LoopBlock.scala 900:55]
  wire  _GEN_163; // @[LoopBlock.scala 900:55]
  wire  _GEN_164; // @[LoopBlock.scala 900:55]
  wire  _GEN_165; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_166; // @[LoopBlock.scala 900:55]
  wire  _GEN_167; // @[LoopBlock.scala 900:55]
  wire  _GEN_168; // @[LoopBlock.scala 900:55]
  wire  _GEN_170; // @[LoopBlock.scala 900:55]
  wire  _GEN_171; // @[LoopBlock.scala 900:55]
  wire [1:0] _GEN_172; // @[LoopBlock.scala 900:55]
  wire  _GEN_173; // @[LoopBlock.scala 900:55]
  wire  _GEN_174; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_175; // @[LoopBlock.scala 900:55]
  wire  _T_830; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_176; // @[LoopBlock.scala 955:48]
  wire  _GEN_177; // @[LoopBlock.scala 955:48]
  wire  _GEN_178; // @[LoopBlock.scala 955:48]
  wire  _GEN_179; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_180; // @[LoopBlock.scala 955:48]
  wire  _GEN_181; // @[LoopBlock.scala 955:48]
  wire  _GEN_182; // @[LoopBlock.scala 955:48]
  wire  _GEN_184; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_185; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_188; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_189; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_191; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_192; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_194; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_197; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_200; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_201; // @[LoopBlock.scala 955:48]
  wire  _GEN_203; // @[LoopBlock.scala 955:48]
  wire  _GEN_204; // @[LoopBlock.scala 955:48]
  wire  _GEN_205; // @[LoopBlock.scala 955:48]
  wire  _GEN_206; // @[LoopBlock.scala 955:48]
  wire  _GEN_207; // @[LoopBlock.scala 955:48]
  wire  _GEN_208; // @[LoopBlock.scala 955:48]
  wire  _GEN_209; // @[LoopBlock.scala 955:48]
  wire [1:0] _GEN_210; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_211; // @[Conditional.scala 39:67]
  wire  _GEN_212; // @[Conditional.scala 39:67]
  wire  _GEN_213; // @[Conditional.scala 39:67]
  wire  _GEN_214; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_215; // @[Conditional.scala 39:67]
  wire  _GEN_216; // @[Conditional.scala 39:67]
  wire  _GEN_217; // @[Conditional.scala 39:67]
  wire  _GEN_219; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_220; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_223; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_224; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_226; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_227; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_229; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_232; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_235; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_236; // @[Conditional.scala 39:67]
  wire  _GEN_238; // @[Conditional.scala 39:67]
  wire  _GEN_239; // @[Conditional.scala 39:67]
  wire  _GEN_240; // @[Conditional.scala 39:67]
  wire  _GEN_241; // @[Conditional.scala 39:67]
  wire  _GEN_242; // @[Conditional.scala 39:67]
  wire  _GEN_243; // @[Conditional.scala 39:67]
  wire  _GEN_244; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_245; // @[Conditional.scala 39:67]
  wire  _GEN_246; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_247; // @[Conditional.scala 39:67]
  wire  _GEN_248; // @[Conditional.scala 39:67]
  wire  _GEN_249; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_250; // @[Conditional.scala 39:67]
  wire  _GEN_251; // @[Conditional.scala 39:67]
  wire  _GEN_252; // @[Conditional.scala 39:67]
  wire  _GEN_253; // @[Conditional.scala 39:67]
  wire  _GEN_254; // @[Conditional.scala 39:67]
  wire  _GEN_255; // @[Conditional.scala 39:67]
  wire  _GEN_256; // @[Conditional.scala 39:67]
  wire  _GEN_257; // @[Conditional.scala 39:67]
  wire  _GEN_258; // @[Conditional.scala 39:67]
  wire  _GEN_259; // @[Conditional.scala 39:67]
  wire  _GEN_261; // @[Conditional.scala 39:67]
  wire  _GEN_262; // @[Conditional.scala 39:67]
  wire  _GEN_263; // @[Conditional.scala 39:67]
  wire  _GEN_264; // @[Conditional.scala 39:67]
  wire  _GEN_265; // @[Conditional.scala 39:67]
  wire  _GEN_266; // @[Conditional.scala 39:67]
  wire  _GEN_267; // @[Conditional.scala 39:67]
  wire  _GEN_268; // @[Conditional.scala 39:67]
  wire  _GEN_269; // @[Conditional.scala 39:67]
  wire  _GEN_270; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_271; // @[Conditional.scala 39:67]
  wire  _GEN_272; // @[Conditional.scala 39:67]
  wire  _GEN_273; // @[Conditional.scala 39:67]
  wire  _GEN_275; // @[Conditional.scala 39:67]
  wire  _GEN_276; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_277; // @[Conditional.scala 39:67]
  wire  _GEN_278; // @[Conditional.scala 39:67]
  wire  _GEN_279; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_280; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_281; // @[Conditional.scala 39:67]
  wire  _GEN_282; // @[Conditional.scala 39:67]
  wire  _GEN_283; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_284; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_287; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_288; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_290; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_291; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_293; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_296; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_299; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_300; // @[Conditional.scala 39:67]
  wire  _GEN_302; // @[Conditional.scala 39:67]
  wire  _GEN_303; // @[Conditional.scala 39:67]
  wire  _GEN_304; // @[Conditional.scala 39:67]
  wire  _GEN_305; // @[Conditional.scala 39:67]
  wire  _GEN_306; // @[Conditional.scala 39:67]
  wire  _GEN_307; // @[Conditional.scala 39:67]
  wire  _GEN_308; // @[Conditional.scala 40:58]
  wire  _GEN_309; // @[Conditional.scala 40:58]
  wire  _GEN_310; // @[Conditional.scala 40:58]
  wire  _GEN_311; // @[Conditional.scala 40:58]
  wire  _GEN_312; // @[Conditional.scala 40:58]
  wire  _GEN_313; // @[Conditional.scala 40:58]
  wire  _GEN_314; // @[Conditional.scala 40:58]
  wire  _GEN_315; // @[Conditional.scala 40:58]
  wire  _GEN_316; // @[Conditional.scala 40:58]
  wire  _GEN_317; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_318; // @[Conditional.scala 40:58]
  wire  _GEN_319; // @[Conditional.scala 40:58]
  wire  _GEN_320; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_321; // @[Conditional.scala 40:58]
  wire  _GEN_322; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_323; // @[Conditional.scala 40:58]
  wire  _GEN_324; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_325; // @[Conditional.scala 40:58]
  wire  _GEN_326; // @[Conditional.scala 40:58]
  wire  _GEN_327; // @[Conditional.scala 40:58]
  wire  _GEN_328; // @[Conditional.scala 40:58]
  wire  _GEN_329; // @[Conditional.scala 40:58]
  wire  _GEN_330; // @[Conditional.scala 40:58]
  wire  _GEN_331; // @[Conditional.scala 40:58]
  wire  _GEN_332; // @[Conditional.scala 40:58]
  wire  _GEN_333; // @[Conditional.scala 40:58]
  wire  _GEN_334; // @[Conditional.scala 40:58]
  wire  _GEN_336; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_337; // @[Conditional.scala 40:58]
  wire  _GEN_338; // @[Conditional.scala 40:58]
  wire  _GEN_339; // @[Conditional.scala 40:58]
  wire  _GEN_341; // @[Conditional.scala 40:58]
  wire  _GEN_342; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_343; // @[Conditional.scala 40:58]
  wire  _GEN_344; // @[Conditional.scala 40:58]
  wire  _GEN_345; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_346; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_349; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_350; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_352; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_353; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_355; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_358; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_361; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_362; // @[Conditional.scala 40:58]
  wire  _GEN_364; // @[Conditional.scala 40:58]
  wire  _GEN_365; // @[Conditional.scala 40:58]
  wire  _GEN_366; // @[Conditional.scala 40:58]
  wire  _GEN_367; // @[Conditional.scala 40:58]
  wire  _GEN_368; // @[Conditional.scala 40:58]
  wire  _GEN_369; // @[Conditional.scala 40:58]
  assign _T_671 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_671 ? io_enable_bits_taskID : enable_R_taskID; // @[LoopBlock.scala 596:26]
  assign _GEN_2 = _T_671 ? io_enable_bits_control : enable_R_control; // @[LoopBlock.scala 596:26]
  assign _GEN_3 = _T_671 ? 1'h1 : enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_674 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_674 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_674 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_674 ? 1'h1 : loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_677 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_677 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_677 ? 1'h1 : loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_680 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_680 ? io_InLiveIn_0_bits_data : in_live_in_R_0_data; // @[LoopBlock.scala 623:33]
  assign _GEN_13 = _T_680 ? 1'h1 : in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_683 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_15 = _T_683 ? io_InLiveIn_1_bits_taskID : in_live_in_R_1_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_16 = _T_683 ? io_InLiveIn_1_bits_data : in_live_in_R_1_data; // @[LoopBlock.scala 623:33]
  assign _GEN_17 = _T_683 ? 1'h1 : in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_686 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_19 = _T_686 ? io_InLiveIn_2_bits_taskID : in_live_in_R_2_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_20 = _T_686 ? io_InLiveIn_2_bits_data : in_live_in_R_2_data; // @[LoopBlock.scala 623:33]
  assign _GEN_21 = _T_686 ? 1'h1 : in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_689 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_24 = _T_689 ? io_InLiveIn_3_bits_data : in_live_in_R_3_data; // @[LoopBlock.scala 623:33]
  assign _GEN_25 = _T_689 ? 1'h1 : in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_692 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_28 = _T_692 ? io_InLiveIn_4_bits_data : in_live_in_R_4_data; // @[LoopBlock.scala 623:33]
  assign _GEN_29 = _T_692 ? 1'h1 : in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_695 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 37:37]
  assign _GEN_31 = _T_695 ? io_InLiveIn_5_bits_taskID : in_live_in_R_5_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_32 = _T_695 ? io_InLiveIn_5_bits_data : in_live_in_R_5_data; // @[LoopBlock.scala 623:33]
  assign _GEN_33 = _T_695 ? 1'h1 : in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_698 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_35 = _T_698 ? io_CarryDepenIn_0_bits_taskID : in_carry_in_R_0_taskID; // @[LoopBlock.scala 641:37]
  assign _GEN_36 = _T_698 ? io_CarryDepenIn_0_bits_data : in_carry_in_R_0_data; // @[LoopBlock.scala 641:37]
  assign _GEN_37 = _T_698 ? 1'h1 : in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_700 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 37:37]
  assign _GEN_38 = _T_700 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_702 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 37:37]
  assign _GEN_39 = _T_702 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_704 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_40 = _T_704 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_41 = _T_704 ? 1'h1 : loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_707 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_42 = _T_707 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_43 = _T_707 ? 1'h1 : out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_710 = io_OutLiveIn_field0_1_ready & io_OutLiveIn_field0_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_44 = _T_710 ? 1'h0 : out_live_in_valid_R_0_1; // @[LoopBlock.scala 722:57]
  assign _GEN_45 = _T_710 ? 1'h1 : out_live_in_fire_R_0_1; // @[LoopBlock.scala 722:57]
  assign _T_713 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_46 = _T_713 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_47 = _T_713 ? 1'h1 : out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_716 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_48 = _T_716 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_49 = _T_716 ? 1'h1 : out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_719 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_50 = _T_719 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_51 = _T_719 ? 1'h1 : out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_722 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_52 = _T_722 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_53 = _T_722 ? 1'h1 : out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_725 = io_OutLiveIn_field4_1_ready & io_OutLiveIn_field4_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_54 = _T_725 ? 1'h0 : out_live_in_valid_R_4_1; // @[LoopBlock.scala 722:57]
  assign _GEN_55 = _T_725 ? 1'h1 : out_live_in_fire_R_4_1; // @[LoopBlock.scala 722:57]
  assign _T_728 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_56 = _T_728 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_57 = _T_728 ? 1'h1 : out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_731 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_58 = _T_731 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_735 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_736 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_737 = _T_736 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_738 = _T_737 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_739 = _T_738 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_740 = _T_739 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_741 = _T_740 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_60 = enable_R_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_61 = enable_R_control ? 1'h1 : _GEN_44; // @[LoopBlock.scala 870:26]
  assign _GEN_62 = enable_R_control ? 1'h1 : _GEN_46; // @[LoopBlock.scala 870:26]
  assign _GEN_63 = enable_R_control ? 1'h1 : _GEN_48; // @[LoopBlock.scala 870:26]
  assign _GEN_64 = enable_R_control ? 1'h1 : _GEN_50; // @[LoopBlock.scala 870:26]
  assign _GEN_65 = enable_R_control ? 1'h1 : _GEN_52; // @[LoopBlock.scala 870:26]
  assign _GEN_66 = enable_R_control ? 1'h1 : _GEN_54; // @[LoopBlock.scala 870:26]
  assign _GEN_67 = enable_R_control ? 1'h1 : _GEN_56; // @[LoopBlock.scala 870:26]
  assign _GEN_68 = enable_R_control ? 1'h1 : _GEN_58; // @[LoopBlock.scala 870:26]
  assign _GEN_69 = enable_R_control ? 1'h1 : active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_70 = enable_R_control ? enable_R_taskID : active_loop_start_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_71 = enable_R_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_72 = enable_R_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_73 = enable_R_control ? enable_R_taskID : active_loop_back_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_74 = enable_R_control ? 1'h1 : _GEN_39; // @[LoopBlock.scala 870:26]
  assign _GEN_75 = enable_R_control ? 2'h1 : 2'h2; // @[LoopBlock.scala 870:26]
  assign _GEN_76 = enable_R_control ? loop_exit_R_0_control : 1'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_77 = enable_R_control ? loop_exit_R_0_taskID : 10'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_78 = enable_R_control ? _GEN_40 : 1'h1; // @[LoopBlock.scala 870:26]
  assign _GEN_79 = _T_741 ? _GEN_60 : _GEN_42; // @[LoopBlock.scala 869:48]
  assign _GEN_80 = _T_741 ? _GEN_61 : _GEN_44; // @[LoopBlock.scala 869:48]
  assign _GEN_81 = _T_741 ? _GEN_62 : _GEN_46; // @[LoopBlock.scala 869:48]
  assign _GEN_82 = _T_741 ? _GEN_63 : _GEN_48; // @[LoopBlock.scala 869:48]
  assign _GEN_83 = _T_741 ? _GEN_64 : _GEN_50; // @[LoopBlock.scala 869:48]
  assign _GEN_84 = _T_741 ? _GEN_65 : _GEN_52; // @[LoopBlock.scala 869:48]
  assign _GEN_85 = _T_741 ? _GEN_66 : _GEN_54; // @[LoopBlock.scala 869:48]
  assign _GEN_86 = _T_741 ? _GEN_67 : _GEN_56; // @[LoopBlock.scala 869:48]
  assign _GEN_87 = _T_741 ? _GEN_68 : _GEN_58; // @[LoopBlock.scala 869:48]
  assign _GEN_88 = _T_741 ? _GEN_69 : active_loop_start_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_89 = _T_741 ? _GEN_70 : active_loop_start_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_90 = _T_741 ? _GEN_71 : _GEN_38; // @[LoopBlock.scala 869:48]
  assign _GEN_91 = _T_741 ? _GEN_72 : active_loop_back_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_92 = _T_741 ? _GEN_73 : active_loop_back_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_93 = _T_741 ? _GEN_74 : _GEN_39; // @[LoopBlock.scala 869:48]
  assign _GEN_94 = _T_741 ? _GEN_75 : state; // @[LoopBlock.scala 869:48]
  assign _GEN_95 = _T_741 ? _GEN_76 : loop_exit_R_0_control; // @[LoopBlock.scala 869:48]
  assign _GEN_96 = _T_741 ? _GEN_77 : loop_exit_R_0_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_97 = _T_741 ? _GEN_78 : _GEN_40; // @[LoopBlock.scala 869:48]
  assign _T_764 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_765 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_768 = out_live_in_fire_R_0_0 & out_live_in_fire_R_0_1; // @[LoopBlock.scala 825:65]
  assign _T_769 = out_live_in_fire_R_4_0 & out_live_in_fire_R_4_1; // @[LoopBlock.scala 825:65]
  assign _T_770 = _T_768 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_771 = _T_770 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_772 = _T_771 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_773 = _T_772 & _T_769; // @[LoopBlock.scala 828:26]
  assign _T_774 = _T_773 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_775 = _T_765 & _T_774; // @[LoopBlock.scala 899:29]
  assign _GEN_98 = loop_finish_R_0_control ? 1'h1 : _GEN_40; // @[LoopBlock.scala 936:64]
  assign _GEN_99 = loop_finish_R_0_control ? 1'h0 : active_loop_start_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_100 = loop_finish_R_0_control ? 10'h0 : active_loop_start_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_101 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_102 = loop_finish_R_0_control ? 10'h0 : active_loop_back_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_103 = loop_finish_R_0_control ? 1'h1 : loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_104 = loop_finish_R_0_control ? loop_back_R_0_taskID : loop_exit_R_0_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_105 = loop_finish_R_0_control ? 2'h2 : state; // @[LoopBlock.scala 936:64]
  assign _GEN_106 = loop_back_R_0_control ? 1'h0 : _GEN_99; // @[LoopBlock.scala 903:56]
  assign _GEN_107 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_100; // @[LoopBlock.scala 903:56]
  assign _GEN_108 = loop_back_R_0_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_109 = loop_back_R_0_control ? 1'h1 : _GEN_101; // @[LoopBlock.scala 903:56]
  assign _GEN_110 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_102; // @[LoopBlock.scala 903:56]
  assign _GEN_111 = loop_back_R_0_control ? 1'h1 : _GEN_39; // @[LoopBlock.scala 903:56]
  assign _GEN_112 = loop_back_R_0_control ? 1'h0 : _GEN_43; // @[LoopBlock.scala 903:56]
  assign _GEN_113 = loop_back_R_0_control ? 1'h0 : _GEN_45; // @[LoopBlock.scala 903:56]
  assign _GEN_114 = loop_back_R_0_control ? 1'h0 : _GEN_47; // @[LoopBlock.scala 903:56]
  assign _GEN_115 = loop_back_R_0_control ? 1'h0 : _GEN_49; // @[LoopBlock.scala 903:56]
  assign _GEN_116 = loop_back_R_0_control ? 1'h0 : _GEN_51; // @[LoopBlock.scala 903:56]
  assign _GEN_117 = loop_back_R_0_control ? 1'h0 : _GEN_53; // @[LoopBlock.scala 903:56]
  assign _GEN_118 = loop_back_R_0_control ? 1'h0 : _GEN_55; // @[LoopBlock.scala 903:56]
  assign _GEN_119 = loop_back_R_0_control ? 1'h0 : _GEN_57; // @[LoopBlock.scala 903:56]
  assign _GEN_121 = loop_back_R_0_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_122 = loop_back_R_0_control ? 1'h1 : _GEN_44; // @[LoopBlock.scala 903:56]
  assign _GEN_123 = loop_back_R_0_control ? 1'h1 : _GEN_46; // @[LoopBlock.scala 903:56]
  assign _GEN_124 = loop_back_R_0_control ? 1'h1 : _GEN_48; // @[LoopBlock.scala 903:56]
  assign _GEN_125 = loop_back_R_0_control ? 1'h1 : _GEN_50; // @[LoopBlock.scala 903:56]
  assign _GEN_126 = loop_back_R_0_control ? 1'h1 : _GEN_52; // @[LoopBlock.scala 903:56]
  assign _GEN_127 = loop_back_R_0_control ? 1'h1 : _GEN_54; // @[LoopBlock.scala 903:56]
  assign _GEN_128 = loop_back_R_0_control ? 1'h1 : _GEN_56; // @[LoopBlock.scala 903:56]
  assign _GEN_129 = loop_back_R_0_control ? 1'h1 : _GEN_58; // @[LoopBlock.scala 903:56]
  assign _GEN_130 = loop_back_R_0_control ? 1'h0 : _GEN_5; // @[LoopBlock.scala 903:56]
  assign _GEN_131 = loop_back_R_0_control ? 10'h0 : _GEN_4; // @[LoopBlock.scala 903:56]
  assign _GEN_132 = loop_back_R_0_control ? 1'h0 : _GEN_6; // @[LoopBlock.scala 903:56]
  assign _GEN_133 = loop_back_R_0_control ? 1'h0 : _GEN_8; // @[LoopBlock.scala 903:56]
  assign _GEN_135 = loop_back_R_0_control ? 1'h0 : _GEN_9; // @[LoopBlock.scala 903:56]
  assign _GEN_136 = loop_back_R_0_control ? 1'h0 : _GEN_37; // @[LoopBlock.scala 903:56]
  assign _GEN_137 = loop_back_R_0_control ? 2'h1 : _GEN_105; // @[LoopBlock.scala 903:56]
  assign _GEN_138 = loop_back_R_0_control ? _GEN_40 : _GEN_98; // @[LoopBlock.scala 903:56]
  assign _GEN_139 = loop_back_R_0_control ? loop_exit_R_0_control : _GEN_103; // @[LoopBlock.scala 903:56]
  assign _GEN_140 = loop_back_R_0_control ? loop_exit_R_0_taskID : _GEN_104; // @[LoopBlock.scala 903:56]
  assign _GEN_141 = _T_775 ? _GEN_106 : active_loop_start_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_142 = _T_775 ? _GEN_107 : active_loop_start_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_143 = _T_775 ? _GEN_108 : _GEN_38; // @[LoopBlock.scala 900:55]
  assign _GEN_144 = _T_775 ? _GEN_109 : active_loop_back_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_145 = _T_775 ? _GEN_110 : active_loop_back_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_146 = _T_775 ? _GEN_111 : _GEN_39; // @[LoopBlock.scala 900:55]
  assign _GEN_147 = _T_775 ? _GEN_112 : _GEN_43; // @[LoopBlock.scala 900:55]
  assign _GEN_148 = _T_775 ? _GEN_113 : _GEN_45; // @[LoopBlock.scala 900:55]
  assign _GEN_149 = _T_775 ? _GEN_114 : _GEN_47; // @[LoopBlock.scala 900:55]
  assign _GEN_150 = _T_775 ? _GEN_115 : _GEN_49; // @[LoopBlock.scala 900:55]
  assign _GEN_151 = _T_775 ? _GEN_116 : _GEN_51; // @[LoopBlock.scala 900:55]
  assign _GEN_152 = _T_775 ? _GEN_117 : _GEN_53; // @[LoopBlock.scala 900:55]
  assign _GEN_153 = _T_775 ? _GEN_118 : _GEN_55; // @[LoopBlock.scala 900:55]
  assign _GEN_154 = _T_775 ? _GEN_119 : _GEN_57; // @[LoopBlock.scala 900:55]
  assign _GEN_156 = _T_775 ? _GEN_121 : _GEN_42; // @[LoopBlock.scala 900:55]
  assign _GEN_157 = _T_775 ? _GEN_122 : _GEN_44; // @[LoopBlock.scala 900:55]
  assign _GEN_158 = _T_775 ? _GEN_123 : _GEN_46; // @[LoopBlock.scala 900:55]
  assign _GEN_159 = _T_775 ? _GEN_124 : _GEN_48; // @[LoopBlock.scala 900:55]
  assign _GEN_160 = _T_775 ? _GEN_125 : _GEN_50; // @[LoopBlock.scala 900:55]
  assign _GEN_161 = _T_775 ? _GEN_126 : _GEN_52; // @[LoopBlock.scala 900:55]
  assign _GEN_162 = _T_775 ? _GEN_127 : _GEN_54; // @[LoopBlock.scala 900:55]
  assign _GEN_163 = _T_775 ? _GEN_128 : _GEN_56; // @[LoopBlock.scala 900:55]
  assign _GEN_164 = _T_775 ? _GEN_129 : _GEN_58; // @[LoopBlock.scala 900:55]
  assign _GEN_165 = _T_775 ? _GEN_130 : _GEN_5; // @[LoopBlock.scala 900:55]
  assign _GEN_166 = _T_775 ? _GEN_131 : _GEN_4; // @[LoopBlock.scala 900:55]
  assign _GEN_167 = _T_775 ? _GEN_132 : _GEN_6; // @[LoopBlock.scala 900:55]
  assign _GEN_168 = _T_775 ? _GEN_133 : _GEN_8; // @[LoopBlock.scala 900:55]
  assign _GEN_170 = _T_775 ? _GEN_135 : _GEN_9; // @[LoopBlock.scala 900:55]
  assign _GEN_171 = _T_775 ? _GEN_136 : _GEN_37; // @[LoopBlock.scala 900:55]
  assign _GEN_172 = _T_775 ? _GEN_137 : state; // @[LoopBlock.scala 900:55]
  assign _GEN_173 = _T_775 ? _GEN_138 : _GEN_40; // @[LoopBlock.scala 900:55]
  assign _GEN_174 = _T_775 ? _GEN_139 : loop_exit_R_0_control; // @[LoopBlock.scala 900:55]
  assign _GEN_175 = _T_775 ? _GEN_140 : loop_exit_R_0_taskID; // @[LoopBlock.scala 900:55]
  assign _T_830 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_176 = loop_exit_fire_R_0 ? 10'h0 : _GEN_1; // @[LoopBlock.scala 955:48]
  assign _GEN_177 = loop_exit_fire_R_0 ? 1'h0 : _GEN_2; // @[LoopBlock.scala 955:48]
  assign _GEN_178 = loop_exit_fire_R_0 ? 1'h0 : _GEN_3; // @[LoopBlock.scala 955:48]
  assign _GEN_179 = loop_exit_fire_R_0 ? 1'h0 : _GEN_5; // @[LoopBlock.scala 955:48]
  assign _GEN_180 = loop_exit_fire_R_0 ? 10'h0 : _GEN_4; // @[LoopBlock.scala 955:48]
  assign _GEN_181 = loop_exit_fire_R_0 ? 1'h0 : _GEN_6; // @[LoopBlock.scala 955:48]
  assign _GEN_182 = loop_exit_fire_R_0 ? 1'h0 : _GEN_8; // @[LoopBlock.scala 955:48]
  assign _GEN_184 = loop_exit_fire_R_0 ? 1'h0 : _GEN_9; // @[LoopBlock.scala 955:48]
  assign _GEN_185 = loop_exit_fire_R_0 ? 32'h0 : _GEN_12; // @[LoopBlock.scala 955:48]
  assign _GEN_188 = loop_exit_fire_R_0 ? 32'h0 : _GEN_16; // @[LoopBlock.scala 955:48]
  assign _GEN_189 = loop_exit_fire_R_0 ? 10'h0 : _GEN_15; // @[LoopBlock.scala 955:48]
  assign _GEN_191 = loop_exit_fire_R_0 ? 32'h0 : _GEN_20; // @[LoopBlock.scala 955:48]
  assign _GEN_192 = loop_exit_fire_R_0 ? 10'h0 : _GEN_19; // @[LoopBlock.scala 955:48]
  assign _GEN_194 = loop_exit_fire_R_0 ? 32'h0 : _GEN_24; // @[LoopBlock.scala 955:48]
  assign _GEN_197 = loop_exit_fire_R_0 ? 32'h0 : _GEN_28; // @[LoopBlock.scala 955:48]
  assign _GEN_200 = loop_exit_fire_R_0 ? 32'h0 : _GEN_32; // @[LoopBlock.scala 955:48]
  assign _GEN_201 = loop_exit_fire_R_0 ? 10'h0 : _GEN_31; // @[LoopBlock.scala 955:48]
  assign _GEN_203 = loop_exit_fire_R_0 ? 1'h0 : _GEN_13; // @[LoopBlock.scala 955:48]
  assign _GEN_204 = loop_exit_fire_R_0 ? 1'h0 : _GEN_17; // @[LoopBlock.scala 955:48]
  assign _GEN_205 = loop_exit_fire_R_0 ? 1'h0 : _GEN_21; // @[LoopBlock.scala 955:48]
  assign _GEN_206 = loop_exit_fire_R_0 ? 1'h0 : _GEN_25; // @[LoopBlock.scala 955:48]
  assign _GEN_207 = loop_exit_fire_R_0 ? 1'h0 : _GEN_29; // @[LoopBlock.scala 955:48]
  assign _GEN_208 = loop_exit_fire_R_0 ? 1'h0 : _GEN_33; // @[LoopBlock.scala 955:48]
  assign _GEN_209 = loop_exit_fire_R_0 ? 1'h0 : _GEN_37; // @[LoopBlock.scala 955:48]
  assign _GEN_210 = loop_exit_fire_R_0 ? 2'h0 : state; // @[LoopBlock.scala 955:48]
  assign _GEN_211 = _T_830 ? _GEN_176 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_212 = _T_830 ? _GEN_177 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_213 = _T_830 ? _GEN_178 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_214 = _T_830 ? _GEN_179 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_215 = _T_830 ? _GEN_180 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_216 = _T_830 ? _GEN_181 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_217 = _T_830 ? _GEN_182 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_219 = _T_830 ? _GEN_184 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_220 = _T_830 ? _GEN_185 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_223 = _T_830 ? _GEN_188 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_224 = _T_830 ? _GEN_189 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_226 = _T_830 ? _GEN_191 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_227 = _T_830 ? _GEN_192 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_229 = _T_830 ? _GEN_194 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_232 = _T_830 ? _GEN_197 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_235 = _T_830 ? _GEN_200 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_236 = _T_830 ? _GEN_201 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_238 = _T_830 ? _GEN_203 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_239 = _T_830 ? _GEN_204 : _GEN_17; // @[Conditional.scala 39:67]
  assign _GEN_240 = _T_830 ? _GEN_205 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_241 = _T_830 ? _GEN_206 : _GEN_25; // @[Conditional.scala 39:67]
  assign _GEN_242 = _T_830 ? _GEN_207 : _GEN_29; // @[Conditional.scala 39:67]
  assign _GEN_243 = _T_830 ? _GEN_208 : _GEN_33; // @[Conditional.scala 39:67]
  assign _GEN_244 = _T_830 ? _GEN_209 : _GEN_37; // @[Conditional.scala 39:67]
  assign _GEN_245 = _T_830 ? _GEN_210 : state; // @[Conditional.scala 39:67]
  assign _GEN_246 = _T_764 ? _GEN_141 : active_loop_start_R_control; // @[Conditional.scala 39:67]
  assign _GEN_247 = _T_764 ? _GEN_142 : active_loop_start_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_248 = _T_764 ? _GEN_143 : _GEN_38; // @[Conditional.scala 39:67]
  assign _GEN_249 = _T_764 ? _GEN_144 : active_loop_back_R_control; // @[Conditional.scala 39:67]
  assign _GEN_250 = _T_764 ? _GEN_145 : active_loop_back_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_251 = _T_764 ? _GEN_146 : _GEN_39; // @[Conditional.scala 39:67]
  assign _GEN_252 = _T_764 ? _GEN_147 : _GEN_43; // @[Conditional.scala 39:67]
  assign _GEN_253 = _T_764 ? _GEN_148 : _GEN_45; // @[Conditional.scala 39:67]
  assign _GEN_254 = _T_764 ? _GEN_149 : _GEN_47; // @[Conditional.scala 39:67]
  assign _GEN_255 = _T_764 ? _GEN_150 : _GEN_49; // @[Conditional.scala 39:67]
  assign _GEN_256 = _T_764 ? _GEN_151 : _GEN_51; // @[Conditional.scala 39:67]
  assign _GEN_257 = _T_764 ? _GEN_152 : _GEN_53; // @[Conditional.scala 39:67]
  assign _GEN_258 = _T_764 ? _GEN_153 : _GEN_55; // @[Conditional.scala 39:67]
  assign _GEN_259 = _T_764 ? _GEN_154 : _GEN_57; // @[Conditional.scala 39:67]
  assign _GEN_261 = _T_764 ? _GEN_156 : _GEN_42; // @[Conditional.scala 39:67]
  assign _GEN_262 = _T_764 ? _GEN_157 : _GEN_44; // @[Conditional.scala 39:67]
  assign _GEN_263 = _T_764 ? _GEN_158 : _GEN_46; // @[Conditional.scala 39:67]
  assign _GEN_264 = _T_764 ? _GEN_159 : _GEN_48; // @[Conditional.scala 39:67]
  assign _GEN_265 = _T_764 ? _GEN_160 : _GEN_50; // @[Conditional.scala 39:67]
  assign _GEN_266 = _T_764 ? _GEN_161 : _GEN_52; // @[Conditional.scala 39:67]
  assign _GEN_267 = _T_764 ? _GEN_162 : _GEN_54; // @[Conditional.scala 39:67]
  assign _GEN_268 = _T_764 ? _GEN_163 : _GEN_56; // @[Conditional.scala 39:67]
  assign _GEN_269 = _T_764 ? _GEN_164 : _GEN_58; // @[Conditional.scala 39:67]
  assign _GEN_270 = _T_764 ? _GEN_165 : _GEN_214; // @[Conditional.scala 39:67]
  assign _GEN_271 = _T_764 ? _GEN_166 : _GEN_215; // @[Conditional.scala 39:67]
  assign _GEN_272 = _T_764 ? _GEN_167 : _GEN_216; // @[Conditional.scala 39:67]
  assign _GEN_273 = _T_764 ? _GEN_168 : _GEN_217; // @[Conditional.scala 39:67]
  assign _GEN_275 = _T_764 ? _GEN_170 : _GEN_219; // @[Conditional.scala 39:67]
  assign _GEN_276 = _T_764 ? _GEN_171 : _GEN_244; // @[Conditional.scala 39:67]
  assign _GEN_277 = _T_764 ? _GEN_172 : _GEN_245; // @[Conditional.scala 39:67]
  assign _GEN_278 = _T_764 ? _GEN_173 : _GEN_40; // @[Conditional.scala 39:67]
  assign _GEN_279 = _T_764 ? _GEN_174 : loop_exit_R_0_control; // @[Conditional.scala 39:67]
  assign _GEN_280 = _T_764 ? _GEN_175 : loop_exit_R_0_taskID; // @[Conditional.scala 39:67]
  assign _GEN_281 = _T_764 ? _GEN_1 : _GEN_211; // @[Conditional.scala 39:67]
  assign _GEN_282 = _T_764 ? _GEN_2 : _GEN_212; // @[Conditional.scala 39:67]
  assign _GEN_283 = _T_764 ? _GEN_3 : _GEN_213; // @[Conditional.scala 39:67]
  assign _GEN_284 = _T_764 ? _GEN_12 : _GEN_220; // @[Conditional.scala 39:67]
  assign _GEN_287 = _T_764 ? _GEN_16 : _GEN_223; // @[Conditional.scala 39:67]
  assign _GEN_288 = _T_764 ? _GEN_15 : _GEN_224; // @[Conditional.scala 39:67]
  assign _GEN_290 = _T_764 ? _GEN_20 : _GEN_226; // @[Conditional.scala 39:67]
  assign _GEN_291 = _T_764 ? _GEN_19 : _GEN_227; // @[Conditional.scala 39:67]
  assign _GEN_293 = _T_764 ? _GEN_24 : _GEN_229; // @[Conditional.scala 39:67]
  assign _GEN_296 = _T_764 ? _GEN_28 : _GEN_232; // @[Conditional.scala 39:67]
  assign _GEN_299 = _T_764 ? _GEN_32 : _GEN_235; // @[Conditional.scala 39:67]
  assign _GEN_300 = _T_764 ? _GEN_31 : _GEN_236; // @[Conditional.scala 39:67]
  assign _GEN_302 = _T_764 ? _GEN_13 : _GEN_238; // @[Conditional.scala 39:67]
  assign _GEN_303 = _T_764 ? _GEN_17 : _GEN_239; // @[Conditional.scala 39:67]
  assign _GEN_304 = _T_764 ? _GEN_21 : _GEN_240; // @[Conditional.scala 39:67]
  assign _GEN_305 = _T_764 ? _GEN_25 : _GEN_241; // @[Conditional.scala 39:67]
  assign _GEN_306 = _T_764 ? _GEN_29 : _GEN_242; // @[Conditional.scala 39:67]
  assign _GEN_307 = _T_764 ? _GEN_33 : _GEN_243; // @[Conditional.scala 39:67]
  assign _GEN_308 = _T_735 ? _GEN_79 : _GEN_261; // @[Conditional.scala 40:58]
  assign _GEN_309 = _T_735 ? _GEN_80 : _GEN_262; // @[Conditional.scala 40:58]
  assign _GEN_310 = _T_735 ? _GEN_81 : _GEN_263; // @[Conditional.scala 40:58]
  assign _GEN_311 = _T_735 ? _GEN_82 : _GEN_264; // @[Conditional.scala 40:58]
  assign _GEN_312 = _T_735 ? _GEN_83 : _GEN_265; // @[Conditional.scala 40:58]
  assign _GEN_313 = _T_735 ? _GEN_84 : _GEN_266; // @[Conditional.scala 40:58]
  assign _GEN_314 = _T_735 ? _GEN_85 : _GEN_267; // @[Conditional.scala 40:58]
  assign _GEN_315 = _T_735 ? _GEN_86 : _GEN_268; // @[Conditional.scala 40:58]
  assign _GEN_316 = _T_735 ? _GEN_87 : _GEN_269; // @[Conditional.scala 40:58]
  assign _GEN_317 = _T_735 ? _GEN_88 : _GEN_246; // @[Conditional.scala 40:58]
  assign _GEN_318 = _T_735 ? _GEN_89 : _GEN_247; // @[Conditional.scala 40:58]
  assign _GEN_319 = _T_735 ? _GEN_90 : _GEN_248; // @[Conditional.scala 40:58]
  assign _GEN_320 = _T_735 ? _GEN_91 : _GEN_249; // @[Conditional.scala 40:58]
  assign _GEN_321 = _T_735 ? _GEN_92 : _GEN_250; // @[Conditional.scala 40:58]
  assign _GEN_322 = _T_735 ? _GEN_93 : _GEN_251; // @[Conditional.scala 40:58]
  assign _GEN_323 = _T_735 ? _GEN_94 : _GEN_277; // @[Conditional.scala 40:58]
  assign _GEN_324 = _T_735 ? _GEN_95 : _GEN_279; // @[Conditional.scala 40:58]
  assign _GEN_325 = _T_735 ? _GEN_96 : _GEN_280; // @[Conditional.scala 40:58]
  assign _GEN_326 = _T_735 ? _GEN_97 : _GEN_278; // @[Conditional.scala 40:58]
  assign _GEN_327 = _T_735 ? _GEN_43 : _GEN_252; // @[Conditional.scala 40:58]
  assign _GEN_328 = _T_735 ? _GEN_45 : _GEN_253; // @[Conditional.scala 40:58]
  assign _GEN_329 = _T_735 ? _GEN_47 : _GEN_254; // @[Conditional.scala 40:58]
  assign _GEN_330 = _T_735 ? _GEN_49 : _GEN_255; // @[Conditional.scala 40:58]
  assign _GEN_331 = _T_735 ? _GEN_51 : _GEN_256; // @[Conditional.scala 40:58]
  assign _GEN_332 = _T_735 ? _GEN_53 : _GEN_257; // @[Conditional.scala 40:58]
  assign _GEN_333 = _T_735 ? _GEN_55 : _GEN_258; // @[Conditional.scala 40:58]
  assign _GEN_334 = _T_735 ? _GEN_57 : _GEN_259; // @[Conditional.scala 40:58]
  assign _GEN_336 = _T_735 ? _GEN_5 : _GEN_270; // @[Conditional.scala 40:58]
  assign _GEN_337 = _T_735 ? _GEN_4 : _GEN_271; // @[Conditional.scala 40:58]
  assign _GEN_338 = _T_735 ? _GEN_6 : _GEN_272; // @[Conditional.scala 40:58]
  assign _GEN_339 = _T_735 ? _GEN_8 : _GEN_273; // @[Conditional.scala 40:58]
  assign _GEN_341 = _T_735 ? _GEN_9 : _GEN_275; // @[Conditional.scala 40:58]
  assign _GEN_342 = _T_735 ? _GEN_37 : _GEN_276; // @[Conditional.scala 40:58]
  assign _GEN_343 = _T_735 ? _GEN_1 : _GEN_281; // @[Conditional.scala 40:58]
  assign _GEN_344 = _T_735 ? _GEN_2 : _GEN_282; // @[Conditional.scala 40:58]
  assign _GEN_345 = _T_735 ? _GEN_3 : _GEN_283; // @[Conditional.scala 40:58]
  assign _GEN_346 = _T_735 ? _GEN_12 : _GEN_284; // @[Conditional.scala 40:58]
  assign _GEN_349 = _T_735 ? _GEN_16 : _GEN_287; // @[Conditional.scala 40:58]
  assign _GEN_350 = _T_735 ? _GEN_15 : _GEN_288; // @[Conditional.scala 40:58]
  assign _GEN_352 = _T_735 ? _GEN_20 : _GEN_290; // @[Conditional.scala 40:58]
  assign _GEN_353 = _T_735 ? _GEN_19 : _GEN_291; // @[Conditional.scala 40:58]
  assign _GEN_355 = _T_735 ? _GEN_24 : _GEN_293; // @[Conditional.scala 40:58]
  assign _GEN_358 = _T_735 ? _GEN_28 : _GEN_296; // @[Conditional.scala 40:58]
  assign _GEN_361 = _T_735 ? _GEN_32 : _GEN_299; // @[Conditional.scala 40:58]
  assign _GEN_362 = _T_735 ? _GEN_31 : _GEN_300; // @[Conditional.scala 40:58]
  assign _GEN_364 = _T_735 ? _GEN_13 : _GEN_302; // @[Conditional.scala 40:58]
  assign _GEN_365 = _T_735 ? _GEN_17 : _GEN_303; // @[Conditional.scala 40:58]
  assign _GEN_366 = _T_735 ? _GEN_21 : _GEN_304; // @[Conditional.scala 40:58]
  assign _GEN_367 = _T_735 ? _GEN_25 : _GEN_305; // @[Conditional.scala 40:58]
  assign _GEN_368 = _T_735 ? _GEN_29 : _GEN_306; // @[Conditional.scala 40:58]
  assign _GEN_369 = _T_735 ? _GEN_33 : _GEN_307; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_taskID = in_live_in_R_5_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_1_valid = out_live_in_valid_R_4_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_1_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_1_valid = out_live_in_valid_R_0_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_1_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_5_taskID = _RAND_15[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_23[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_0_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_live_in_valid_R_4_1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_live_in_fire_R_0_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  out_live_in_fire_R_4_1 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_43[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_46[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_49[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  state = _RAND_53[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_671) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_764) begin
          if (_T_671) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_671) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_671) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_671) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_764) begin
          if (_T_671) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_671) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_671) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_671) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_671) begin
            enable_valid_R <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_671) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_671) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_674) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_674) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_674) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_674) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_674) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_674) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_674) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_674) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_674) begin
          loop_back_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_674) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_674) begin
              loop_back_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_674) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_677) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_677) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_677) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_677) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_8;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_677) begin
          loop_finish_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_677) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_677) begin
              loop_finish_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_677) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_735) begin
        if (_T_680) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_764) begin
          if (_T_680) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_680) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_680) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_683) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_764) begin
          if (_T_683) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_taskID <= 10'h0;
            end else begin
              if (_T_683) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_683) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_735) begin
        if (_T_683) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_764) begin
          if (_T_683) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_683) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_683) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_686) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_764) begin
          if (_T_686) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_taskID <= 10'h0;
            end else begin
              if (_T_686) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_686) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_735) begin
        if (_T_686) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_764) begin
          if (_T_686) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_686) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_686) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_735) begin
        if (_T_689) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_764) begin
          if (_T_689) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_689) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_689) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_735) begin
        if (_T_692) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_764) begin
          if (_T_692) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_692) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_692) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_695) begin
          in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
        end
      end else begin
        if (_T_764) begin
          if (_T_695) begin
            in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_taskID <= 10'h0;
            end else begin
              if (_T_695) begin
                in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
              end
            end
          end else begin
            if (_T_695) begin
              in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_735) begin
        if (_T_695) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_764) begin
          if (_T_695) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_695) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_695) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_680) begin
          in_live_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_680) begin
            in_live_in_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_680) begin
                in_live_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_680) begin
              in_live_in_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_683) begin
          in_live_in_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_683) begin
            in_live_in_valid_R_1 <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              if (_T_683) begin
                in_live_in_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_683) begin
              in_live_in_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_686) begin
          in_live_in_valid_R_2 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_686) begin
            in_live_in_valid_R_2 <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              if (_T_686) begin
                in_live_in_valid_R_2 <= 1'h1;
              end
            end
          end else begin
            if (_T_686) begin
              in_live_in_valid_R_2 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_689) begin
          in_live_in_valid_R_3 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_689) begin
            in_live_in_valid_R_3 <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              if (_T_689) begin
                in_live_in_valid_R_3 <= 1'h1;
              end
            end
          end else begin
            if (_T_689) begin
              in_live_in_valid_R_3 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_692) begin
          in_live_in_valid_R_4 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_692) begin
            in_live_in_valid_R_4 <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              if (_T_692) begin
                in_live_in_valid_R_4 <= 1'h1;
              end
            end
          end else begin
            if (_T_692) begin
              in_live_in_valid_R_4 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_695) begin
          in_live_in_valid_R_5 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_695) begin
            in_live_in_valid_R_5 <= 1'h1;
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              if (_T_695) begin
                in_live_in_valid_R_5 <= 1'h1;
              end
            end
          end else begin
            if (_T_695) begin
              in_live_in_valid_R_5 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_698) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_698) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_698) begin
          in_carry_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_698) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_698) begin
              in_carry_in_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_698) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_707) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_707) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_707) begin
                out_live_in_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_707) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_0_0 <= _GEN_42;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_1 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_0_1 <= 1'h1;
          end else begin
            if (_T_710) begin
              out_live_in_valid_R_0_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_710) begin
            out_live_in_valid_R_0_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_0_1 <= 1'h1;
            end else begin
              if (_T_710) begin
                out_live_in_valid_R_0_1 <= 1'h0;
              end
            end
          end else begin
            if (_T_710) begin
              out_live_in_valid_R_0_1 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_0_1 <= _GEN_44;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_1_0 <= 1'h1;
          end else begin
            if (_T_713) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_713) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_1_0 <= 1'h1;
            end else begin
              if (_T_713) begin
                out_live_in_valid_R_1_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_713) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_1_0 <= _GEN_46;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_2_0 <= 1'h1;
          end else begin
            if (_T_716) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_716) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_2_0 <= 1'h1;
            end else begin
              if (_T_716) begin
                out_live_in_valid_R_2_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_716) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_2_0 <= _GEN_48;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_3_0 <= 1'h1;
          end else begin
            if (_T_719) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_719) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_3_0 <= 1'h1;
            end else begin
              if (_T_719) begin
                out_live_in_valid_R_3_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_719) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_3_0 <= _GEN_50;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_4_0 <= 1'h1;
          end else begin
            if (_T_722) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_722) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_4_0 <= 1'h1;
            end else begin
              if (_T_722) begin
                out_live_in_valid_R_4_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_722) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_4_0 <= _GEN_52;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_1 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_4_1 <= 1'h1;
          end else begin
            if (_T_725) begin
              out_live_in_valid_R_4_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_725) begin
            out_live_in_valid_R_4_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_4_1 <= 1'h1;
            end else begin
              if (_T_725) begin
                out_live_in_valid_R_4_1 <= 1'h0;
              end
            end
          end else begin
            if (_T_725) begin
              out_live_in_valid_R_4_1 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_4_1 <= _GEN_54;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_live_in_valid_R_5_0 <= 1'h1;
          end else begin
            if (_T_728) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_728) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_5_0 <= 1'h1;
            end else begin
              if (_T_728) begin
                out_live_in_valid_R_5_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_728) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_5_0 <= _GEN_56;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_707) begin
          out_live_in_fire_R_0_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              if (_T_707) begin
                out_live_in_fire_R_0_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_707) begin
              out_live_in_fire_R_0_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_707) begin
            out_live_in_fire_R_0_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_1 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_710) begin
          out_live_in_fire_R_0_1 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_1 <= 1'h0;
            end else begin
              if (_T_710) begin
                out_live_in_fire_R_0_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_710) begin
              out_live_in_fire_R_0_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_710) begin
            out_live_in_fire_R_0_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_713) begin
          out_live_in_fire_R_1_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              if (_T_713) begin
                out_live_in_fire_R_1_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_713) begin
              out_live_in_fire_R_1_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_713) begin
            out_live_in_fire_R_1_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_716) begin
          out_live_in_fire_R_2_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              if (_T_716) begin
                out_live_in_fire_R_2_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_716) begin
              out_live_in_fire_R_2_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_716) begin
            out_live_in_fire_R_2_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_719) begin
          out_live_in_fire_R_3_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              if (_T_719) begin
                out_live_in_fire_R_3_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_719) begin
              out_live_in_fire_R_3_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_719) begin
            out_live_in_fire_R_3_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_722) begin
          out_live_in_fire_R_4_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              if (_T_722) begin
                out_live_in_fire_R_4_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_722) begin
              out_live_in_fire_R_4_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_722) begin
            out_live_in_fire_R_4_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_1 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_725) begin
          out_live_in_fire_R_4_1 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_1 <= 1'h0;
            end else begin
              if (_T_725) begin
                out_live_in_fire_R_4_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_725) begin
              out_live_in_fire_R_4_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_725) begin
            out_live_in_fire_R_4_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_728) begin
          out_live_in_fire_R_5_0 <= 1'h1;
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              if (_T_728) begin
                out_live_in_fire_R_5_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_728) begin
              out_live_in_fire_R_5_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_728) begin
            out_live_in_fire_R_5_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            out_carry_out_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_731) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_731) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              out_carry_out_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_731) begin
                out_carry_out_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_731) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_carry_out_valid_R_0_0 <= _GEN_58;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            active_loop_start_R_control <= 1'h1;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            active_loop_start_valid_R <= 1'h1;
          end else begin
            if (_T_700) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_700) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              active_loop_start_valid_R <= 1'h1;
            end else begin
              if (_T_700) begin
                active_loop_start_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_700) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_start_valid_R <= _GEN_38;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_control <= 1'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            active_loop_back_valid_R <= 1'h1;
          end else begin
            if (_T_702) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_702) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              active_loop_back_valid_R <= 1'h1;
            end else begin
              if (_T_702) begin
                active_loop_back_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_702) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_back_valid_R <= _GEN_39;
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 10'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 10'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_control <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_control <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            if (_T_704) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_704) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              if (_T_704) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              if (loop_finish_R_0_control) begin
                loop_exit_valid_R_0 <= 1'h1;
              end else begin
                if (_T_704) begin
                  loop_exit_valid_R_0 <= 1'h0;
                end
              end
            end
          end else begin
            loop_exit_valid_R_0 <= _GEN_40;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      if (_T_704) begin
        loop_exit_fire_R_0 <= 1'h1;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_735) begin
        if (_T_741) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_764) begin
          if (_T_775) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_830) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [9:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [9:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [9:0]  io_InLiveIn_3_bits_taskID,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [31:0] io_InLiveIn_4_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [9:0]  io_OutLiveIn_field3_0_bits_taskID,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [9:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [9:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [9:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [9:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [9:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [9:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [9:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [9:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_2;
  reg [9:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_3;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_5;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_6;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_7;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_8;
  reg [9:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [9:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [9:0] in_live_in_R_3_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_16;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_17;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_18;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_19;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_20;
  reg [9:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_21;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_22;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_23;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_24;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_25;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_26;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_29;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_30;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_31;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_32;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_33;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_34;
  reg [9:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_35;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_36;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_37;
  reg [9:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_38;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_39;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_40;
  reg [9:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_41;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_42;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_43;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_44;
  wire  _T_577; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[LoopBlock.scala 596:26]
  wire  _GEN_2; // @[LoopBlock.scala 596:26]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_580; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_4; // @[LoopBlock.scala 603:33]
  wire  _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_583; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_586; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[LoopBlock.scala 623:33]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_589; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_15; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_16; // @[LoopBlock.scala 623:33]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_592; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_19; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_20; // @[LoopBlock.scala 623:33]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_595; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_23; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_24; // @[LoopBlock.scala 623:33]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_598; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_28; // @[LoopBlock.scala 623:33]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_601; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_31; // @[LoopBlock.scala 641:37]
  wire [31:0] _GEN_32; // @[LoopBlock.scala 641:37]
  wire  _GEN_33; // @[LoopBlock.scala 641:37]
  wire  _T_603; // @[Decoupled.scala 37:37]
  wire  _GEN_34; // @[LoopBlock.scala 704:39]
  wire  _T_605; // @[Decoupled.scala 37:37]
  wire  _GEN_35; // @[LoopBlock.scala 708:38]
  wire  _T_607; // @[Decoupled.scala 37:37]
  wire  _GEN_36; // @[LoopBlock.scala 713:33]
  wire  _GEN_37; // @[LoopBlock.scala 713:33]
  wire  _T_610; // @[Decoupled.scala 37:37]
  wire  _GEN_38; // @[LoopBlock.scala 722:57]
  wire  _GEN_39; // @[LoopBlock.scala 722:57]
  wire  _T_613; // @[Decoupled.scala 37:37]
  wire  _GEN_40; // @[LoopBlock.scala 722:57]
  wire  _GEN_41; // @[LoopBlock.scala 722:57]
  wire  _T_616; // @[Decoupled.scala 37:37]
  wire  _GEN_42; // @[LoopBlock.scala 722:57]
  wire  _GEN_43; // @[LoopBlock.scala 722:57]
  wire  _T_619; // @[Decoupled.scala 37:37]
  wire  _GEN_44; // @[LoopBlock.scala 722:57]
  wire  _GEN_45; // @[LoopBlock.scala 722:57]
  wire  _T_622; // @[Decoupled.scala 37:37]
  wire  _GEN_46; // @[LoopBlock.scala 722:57]
  wire  _GEN_47; // @[LoopBlock.scala 722:57]
  wire  _T_625; // @[Decoupled.scala 37:37]
  wire  _GEN_48; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_45;
  wire  _T_629; // @[Conditional.scala 37:30]
  wire  _T_630; // @[LoopBlock.scala 765:35]
  wire  _T_631; // @[LoopBlock.scala 765:35]
  wire  _T_632; // @[LoopBlock.scala 765:35]
  wire  _T_633; // @[LoopBlock.scala 765:35]
  wire  _T_634; // @[LoopBlock.scala 869:28]
  wire  _GEN_50; // @[LoopBlock.scala 870:26]
  wire  _GEN_51; // @[LoopBlock.scala 870:26]
  wire  _GEN_52; // @[LoopBlock.scala 870:26]
  wire  _GEN_53; // @[LoopBlock.scala 870:26]
  wire  _GEN_54; // @[LoopBlock.scala 870:26]
  wire  _GEN_55; // @[LoopBlock.scala 870:26]
  wire  _GEN_56; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_57; // @[LoopBlock.scala 870:26]
  wire  _GEN_58; // @[LoopBlock.scala 870:26]
  wire  _GEN_59; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_60; // @[LoopBlock.scala 870:26]
  wire  _GEN_61; // @[LoopBlock.scala 870:26]
  wire [1:0] _GEN_62; // @[LoopBlock.scala 870:26]
  wire  _GEN_63; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_64; // @[LoopBlock.scala 870:26]
  wire  _GEN_65; // @[LoopBlock.scala 870:26]
  wire  _GEN_66; // @[LoopBlock.scala 869:48]
  wire  _GEN_67; // @[LoopBlock.scala 869:48]
  wire  _GEN_68; // @[LoopBlock.scala 869:48]
  wire  _GEN_69; // @[LoopBlock.scala 869:48]
  wire  _GEN_70; // @[LoopBlock.scala 869:48]
  wire  _GEN_71; // @[LoopBlock.scala 869:48]
  wire  _GEN_72; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_73; // @[LoopBlock.scala 869:48]
  wire  _GEN_74; // @[LoopBlock.scala 869:48]
  wire  _GEN_75; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_76; // @[LoopBlock.scala 869:48]
  wire  _GEN_77; // @[LoopBlock.scala 869:48]
  wire [1:0] _GEN_78; // @[LoopBlock.scala 869:48]
  wire  _GEN_79; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_80; // @[LoopBlock.scala 869:48]
  wire  _GEN_81; // @[LoopBlock.scala 869:48]
  wire  _T_654; // @[Conditional.scala 37:30]
  wire  _T_655; // @[LoopBlock.scala 898:30]
  wire  _T_658; // @[LoopBlock.scala 828:26]
  wire  _T_659; // @[LoopBlock.scala 828:26]
  wire  _T_660; // @[LoopBlock.scala 828:26]
  wire  _T_661; // @[LoopBlock.scala 828:26]
  wire  _T_662; // @[LoopBlock.scala 899:29]
  wire  _GEN_82; // @[LoopBlock.scala 936:64]
  wire  _GEN_83; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_84; // @[LoopBlock.scala 936:64]
  wire  _GEN_85; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_86; // @[LoopBlock.scala 936:64]
  wire  _GEN_87; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_88; // @[LoopBlock.scala 936:64]
  wire [1:0] _GEN_89; // @[LoopBlock.scala 936:64]
  wire  _GEN_90; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_91; // @[LoopBlock.scala 903:56]
  wire  _GEN_92; // @[LoopBlock.scala 903:56]
  wire  _GEN_93; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_94; // @[LoopBlock.scala 903:56]
  wire  _GEN_95; // @[LoopBlock.scala 903:56]
  wire  _GEN_96; // @[LoopBlock.scala 903:56]
  wire  _GEN_97; // @[LoopBlock.scala 903:56]
  wire  _GEN_98; // @[LoopBlock.scala 903:56]
  wire  _GEN_99; // @[LoopBlock.scala 903:56]
  wire  _GEN_100; // @[LoopBlock.scala 903:56]
  wire  _GEN_102; // @[LoopBlock.scala 903:56]
  wire  _GEN_103; // @[LoopBlock.scala 903:56]
  wire  _GEN_104; // @[LoopBlock.scala 903:56]
  wire  _GEN_105; // @[LoopBlock.scala 903:56]
  wire  _GEN_106; // @[LoopBlock.scala 903:56]
  wire  _GEN_107; // @[LoopBlock.scala 903:56]
  wire  _GEN_108; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_109; // @[LoopBlock.scala 903:56]
  wire  _GEN_110; // @[LoopBlock.scala 903:56]
  wire  _GEN_111; // @[LoopBlock.scala 903:56]
  wire  _GEN_113; // @[LoopBlock.scala 903:56]
  wire  _GEN_114; // @[LoopBlock.scala 903:56]
  wire [1:0] _GEN_115; // @[LoopBlock.scala 903:56]
  wire  _GEN_116; // @[LoopBlock.scala 903:56]
  wire  _GEN_117; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_118; // @[LoopBlock.scala 903:56]
  wire  _GEN_119; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_120; // @[LoopBlock.scala 900:55]
  wire  _GEN_121; // @[LoopBlock.scala 900:55]
  wire  _GEN_122; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_123; // @[LoopBlock.scala 900:55]
  wire  _GEN_124; // @[LoopBlock.scala 900:55]
  wire  _GEN_125; // @[LoopBlock.scala 900:55]
  wire  _GEN_126; // @[LoopBlock.scala 900:55]
  wire  _GEN_127; // @[LoopBlock.scala 900:55]
  wire  _GEN_128; // @[LoopBlock.scala 900:55]
  wire  _GEN_129; // @[LoopBlock.scala 900:55]
  wire  _GEN_131; // @[LoopBlock.scala 900:55]
  wire  _GEN_132; // @[LoopBlock.scala 900:55]
  wire  _GEN_133; // @[LoopBlock.scala 900:55]
  wire  _GEN_134; // @[LoopBlock.scala 900:55]
  wire  _GEN_135; // @[LoopBlock.scala 900:55]
  wire  _GEN_136; // @[LoopBlock.scala 900:55]
  wire  _GEN_137; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_138; // @[LoopBlock.scala 900:55]
  wire  _GEN_139; // @[LoopBlock.scala 900:55]
  wire  _GEN_140; // @[LoopBlock.scala 900:55]
  wire  _GEN_142; // @[LoopBlock.scala 900:55]
  wire  _GEN_143; // @[LoopBlock.scala 900:55]
  wire [1:0] _GEN_144; // @[LoopBlock.scala 900:55]
  wire  _GEN_145; // @[LoopBlock.scala 900:55]
  wire  _GEN_146; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_147; // @[LoopBlock.scala 900:55]
  wire  _T_711; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_148; // @[LoopBlock.scala 955:48]
  wire  _GEN_149; // @[LoopBlock.scala 955:48]
  wire  _GEN_150; // @[LoopBlock.scala 955:48]
  wire  _GEN_151; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_152; // @[LoopBlock.scala 955:48]
  wire  _GEN_153; // @[LoopBlock.scala 955:48]
  wire  _GEN_154; // @[LoopBlock.scala 955:48]
  wire  _GEN_156; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_157; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_160; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_161; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_163; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_164; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_166; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_167; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_169; // @[LoopBlock.scala 955:48]
  wire  _GEN_172; // @[LoopBlock.scala 955:48]
  wire  _GEN_173; // @[LoopBlock.scala 955:48]
  wire  _GEN_174; // @[LoopBlock.scala 955:48]
  wire  _GEN_175; // @[LoopBlock.scala 955:48]
  wire  _GEN_176; // @[LoopBlock.scala 955:48]
  wire  _GEN_177; // @[LoopBlock.scala 955:48]
  wire [1:0] _GEN_178; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_179; // @[Conditional.scala 39:67]
  wire  _GEN_180; // @[Conditional.scala 39:67]
  wire  _GEN_181; // @[Conditional.scala 39:67]
  wire  _GEN_182; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_183; // @[Conditional.scala 39:67]
  wire  _GEN_184; // @[Conditional.scala 39:67]
  wire  _GEN_185; // @[Conditional.scala 39:67]
  wire  _GEN_187; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_188; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_191; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_192; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_194; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_195; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_197; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_198; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_200; // @[Conditional.scala 39:67]
  wire  _GEN_203; // @[Conditional.scala 39:67]
  wire  _GEN_204; // @[Conditional.scala 39:67]
  wire  _GEN_205; // @[Conditional.scala 39:67]
  wire  _GEN_206; // @[Conditional.scala 39:67]
  wire  _GEN_207; // @[Conditional.scala 39:67]
  wire  _GEN_208; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_209; // @[Conditional.scala 39:67]
  wire  _GEN_210; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_211; // @[Conditional.scala 39:67]
  wire  _GEN_212; // @[Conditional.scala 39:67]
  wire  _GEN_213; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_214; // @[Conditional.scala 39:67]
  wire  _GEN_215; // @[Conditional.scala 39:67]
  wire  _GEN_216; // @[Conditional.scala 39:67]
  wire  _GEN_217; // @[Conditional.scala 39:67]
  wire  _GEN_218; // @[Conditional.scala 39:67]
  wire  _GEN_219; // @[Conditional.scala 39:67]
  wire  _GEN_220; // @[Conditional.scala 39:67]
  wire  _GEN_222; // @[Conditional.scala 39:67]
  wire  _GEN_223; // @[Conditional.scala 39:67]
  wire  _GEN_224; // @[Conditional.scala 39:67]
  wire  _GEN_225; // @[Conditional.scala 39:67]
  wire  _GEN_226; // @[Conditional.scala 39:67]
  wire  _GEN_227; // @[Conditional.scala 39:67]
  wire  _GEN_228; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_229; // @[Conditional.scala 39:67]
  wire  _GEN_230; // @[Conditional.scala 39:67]
  wire  _GEN_231; // @[Conditional.scala 39:67]
  wire  _GEN_233; // @[Conditional.scala 39:67]
  wire  _GEN_234; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_235; // @[Conditional.scala 39:67]
  wire  _GEN_236; // @[Conditional.scala 39:67]
  wire  _GEN_237; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_238; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_239; // @[Conditional.scala 39:67]
  wire  _GEN_240; // @[Conditional.scala 39:67]
  wire  _GEN_241; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_242; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_245; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_246; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_248; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_249; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_251; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_252; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_254; // @[Conditional.scala 39:67]
  wire  _GEN_257; // @[Conditional.scala 39:67]
  wire  _GEN_258; // @[Conditional.scala 39:67]
  wire  _GEN_259; // @[Conditional.scala 39:67]
  wire  _GEN_260; // @[Conditional.scala 39:67]
  wire  _GEN_261; // @[Conditional.scala 39:67]
  wire  _GEN_262; // @[Conditional.scala 40:58]
  wire  _GEN_263; // @[Conditional.scala 40:58]
  wire  _GEN_264; // @[Conditional.scala 40:58]
  wire  _GEN_265; // @[Conditional.scala 40:58]
  wire  _GEN_266; // @[Conditional.scala 40:58]
  wire  _GEN_267; // @[Conditional.scala 40:58]
  wire  _GEN_268; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_269; // @[Conditional.scala 40:58]
  wire  _GEN_270; // @[Conditional.scala 40:58]
  wire  _GEN_271; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_272; // @[Conditional.scala 40:58]
  wire  _GEN_273; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_274; // @[Conditional.scala 40:58]
  wire  _GEN_275; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_276; // @[Conditional.scala 40:58]
  wire  _GEN_277; // @[Conditional.scala 40:58]
  wire  _GEN_278; // @[Conditional.scala 40:58]
  wire  _GEN_279; // @[Conditional.scala 40:58]
  wire  _GEN_280; // @[Conditional.scala 40:58]
  wire  _GEN_281; // @[Conditional.scala 40:58]
  wire  _GEN_282; // @[Conditional.scala 40:58]
  wire  _GEN_284; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_285; // @[Conditional.scala 40:58]
  wire  _GEN_286; // @[Conditional.scala 40:58]
  wire  _GEN_287; // @[Conditional.scala 40:58]
  wire  _GEN_289; // @[Conditional.scala 40:58]
  wire  _GEN_290; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_291; // @[Conditional.scala 40:58]
  wire  _GEN_292; // @[Conditional.scala 40:58]
  wire  _GEN_293; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_294; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_297; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_298; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_300; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_301; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_303; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_304; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_306; // @[Conditional.scala 40:58]
  wire  _GEN_309; // @[Conditional.scala 40:58]
  wire  _GEN_310; // @[Conditional.scala 40:58]
  wire  _GEN_311; // @[Conditional.scala 40:58]
  wire  _GEN_312; // @[Conditional.scala 40:58]
  wire  _GEN_313; // @[Conditional.scala 40:58]
  assign _T_577 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_577 ? io_enable_bits_taskID : enable_R_taskID; // @[LoopBlock.scala 596:26]
  assign _GEN_2 = _T_577 ? io_enable_bits_control : enable_R_control; // @[LoopBlock.scala 596:26]
  assign _GEN_3 = _T_577 ? 1'h1 : enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_580 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_580 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_580 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_580 ? 1'h1 : loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_583 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_583 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_583 ? 1'h1 : loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_586 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_586 ? io_InLiveIn_0_bits_data : in_live_in_R_0_data; // @[LoopBlock.scala 623:33]
  assign _GEN_13 = _T_586 ? 1'h1 : in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_589 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_15 = _T_589 ? io_InLiveIn_1_bits_taskID : in_live_in_R_1_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_16 = _T_589 ? io_InLiveIn_1_bits_data : in_live_in_R_1_data; // @[LoopBlock.scala 623:33]
  assign _GEN_17 = _T_589 ? 1'h1 : in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_592 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_19 = _T_592 ? io_InLiveIn_2_bits_taskID : in_live_in_R_2_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_20 = _T_592 ? io_InLiveIn_2_bits_data : in_live_in_R_2_data; // @[LoopBlock.scala 623:33]
  assign _GEN_21 = _T_592 ? 1'h1 : in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_595 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_23 = _T_595 ? io_InLiveIn_3_bits_taskID : in_live_in_R_3_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_24 = _T_595 ? io_InLiveIn_3_bits_data : in_live_in_R_3_data; // @[LoopBlock.scala 623:33]
  assign _GEN_25 = _T_595 ? 1'h1 : in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_598 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_28 = _T_598 ? io_InLiveIn_4_bits_data : in_live_in_R_4_data; // @[LoopBlock.scala 623:33]
  assign _GEN_29 = _T_598 ? 1'h1 : in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_601 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_31 = _T_601 ? io_CarryDepenIn_0_bits_taskID : in_carry_in_R_0_taskID; // @[LoopBlock.scala 641:37]
  assign _GEN_32 = _T_601 ? io_CarryDepenIn_0_bits_data : in_carry_in_R_0_data; // @[LoopBlock.scala 641:37]
  assign _GEN_33 = _T_601 ? 1'h1 : in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_603 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 37:37]
  assign _GEN_34 = _T_603 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_605 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 37:37]
  assign _GEN_35 = _T_605 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_607 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_36 = _T_607 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_37 = _T_607 ? 1'h1 : loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_610 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_38 = _T_610 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_39 = _T_610 ? 1'h1 : out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_613 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_40 = _T_613 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_41 = _T_613 ? 1'h1 : out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_616 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_42 = _T_616 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_43 = _T_616 ? 1'h1 : out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_619 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_44 = _T_619 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_45 = _T_619 ? 1'h1 : out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_622 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_46 = _T_622 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_47 = _T_622 ? 1'h1 : out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_625 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_48 = _T_625 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_629 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_630 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_631 = _T_630 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_632 = _T_631 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_633 = _T_632 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_634 = _T_633 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_50 = enable_R_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_51 = enable_R_control ? 1'h1 : _GEN_40; // @[LoopBlock.scala 870:26]
  assign _GEN_52 = enable_R_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_53 = enable_R_control ? 1'h1 : _GEN_44; // @[LoopBlock.scala 870:26]
  assign _GEN_54 = enable_R_control ? 1'h1 : _GEN_46; // @[LoopBlock.scala 870:26]
  assign _GEN_55 = enable_R_control ? 1'h1 : _GEN_48; // @[LoopBlock.scala 870:26]
  assign _GEN_56 = enable_R_control ? 1'h1 : active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_57 = enable_R_control ? enable_R_taskID : active_loop_start_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_58 = enable_R_control ? 1'h1 : _GEN_34; // @[LoopBlock.scala 870:26]
  assign _GEN_59 = enable_R_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_60 = enable_R_control ? enable_R_taskID : active_loop_back_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_61 = enable_R_control ? 1'h1 : _GEN_35; // @[LoopBlock.scala 870:26]
  assign _GEN_62 = enable_R_control ? 2'h1 : 2'h2; // @[LoopBlock.scala 870:26]
  assign _GEN_63 = enable_R_control ? loop_exit_R_0_control : 1'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_64 = enable_R_control ? loop_exit_R_0_taskID : 10'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_65 = enable_R_control ? _GEN_36 : 1'h1; // @[LoopBlock.scala 870:26]
  assign _GEN_66 = _T_634 ? _GEN_50 : _GEN_38; // @[LoopBlock.scala 869:48]
  assign _GEN_67 = _T_634 ? _GEN_51 : _GEN_40; // @[LoopBlock.scala 869:48]
  assign _GEN_68 = _T_634 ? _GEN_52 : _GEN_42; // @[LoopBlock.scala 869:48]
  assign _GEN_69 = _T_634 ? _GEN_53 : _GEN_44; // @[LoopBlock.scala 869:48]
  assign _GEN_70 = _T_634 ? _GEN_54 : _GEN_46; // @[LoopBlock.scala 869:48]
  assign _GEN_71 = _T_634 ? _GEN_55 : _GEN_48; // @[LoopBlock.scala 869:48]
  assign _GEN_72 = _T_634 ? _GEN_56 : active_loop_start_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_73 = _T_634 ? _GEN_57 : active_loop_start_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_74 = _T_634 ? _GEN_58 : _GEN_34; // @[LoopBlock.scala 869:48]
  assign _GEN_75 = _T_634 ? _GEN_59 : active_loop_back_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_76 = _T_634 ? _GEN_60 : active_loop_back_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_77 = _T_634 ? _GEN_61 : _GEN_35; // @[LoopBlock.scala 869:48]
  assign _GEN_78 = _T_634 ? _GEN_62 : state; // @[LoopBlock.scala 869:48]
  assign _GEN_79 = _T_634 ? _GEN_63 : loop_exit_R_0_control; // @[LoopBlock.scala 869:48]
  assign _GEN_80 = _T_634 ? _GEN_64 : loop_exit_R_0_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_81 = _T_634 ? _GEN_65 : _GEN_36; // @[LoopBlock.scala 869:48]
  assign _T_654 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_655 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_658 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_659 = _T_658 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_660 = _T_659 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_661 = _T_660 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_662 = _T_655 & _T_661; // @[LoopBlock.scala 899:29]
  assign _GEN_82 = loop_finish_R_0_control ? 1'h1 : _GEN_36; // @[LoopBlock.scala 936:64]
  assign _GEN_83 = loop_finish_R_0_control ? 1'h0 : active_loop_start_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_84 = loop_finish_R_0_control ? 10'h0 : active_loop_start_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_85 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_86 = loop_finish_R_0_control ? 10'h0 : active_loop_back_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_87 = loop_finish_R_0_control ? 1'h1 : loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_88 = loop_finish_R_0_control ? loop_back_R_0_taskID : loop_exit_R_0_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_89 = loop_finish_R_0_control ? 2'h2 : state; // @[LoopBlock.scala 936:64]
  assign _GEN_90 = loop_back_R_0_control ? 1'h0 : _GEN_83; // @[LoopBlock.scala 903:56]
  assign _GEN_91 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_84; // @[LoopBlock.scala 903:56]
  assign _GEN_92 = loop_back_R_0_control ? 1'h1 : _GEN_34; // @[LoopBlock.scala 903:56]
  assign _GEN_93 = loop_back_R_0_control ? 1'h1 : _GEN_85; // @[LoopBlock.scala 903:56]
  assign _GEN_94 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_86; // @[LoopBlock.scala 903:56]
  assign _GEN_95 = loop_back_R_0_control ? 1'h1 : _GEN_35; // @[LoopBlock.scala 903:56]
  assign _GEN_96 = loop_back_R_0_control ? 1'h0 : _GEN_39; // @[LoopBlock.scala 903:56]
  assign _GEN_97 = loop_back_R_0_control ? 1'h0 : _GEN_41; // @[LoopBlock.scala 903:56]
  assign _GEN_98 = loop_back_R_0_control ? 1'h0 : _GEN_43; // @[LoopBlock.scala 903:56]
  assign _GEN_99 = loop_back_R_0_control ? 1'h0 : _GEN_45; // @[LoopBlock.scala 903:56]
  assign _GEN_100 = loop_back_R_0_control ? 1'h0 : _GEN_47; // @[LoopBlock.scala 903:56]
  assign _GEN_102 = loop_back_R_0_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_103 = loop_back_R_0_control ? 1'h1 : _GEN_40; // @[LoopBlock.scala 903:56]
  assign _GEN_104 = loop_back_R_0_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_105 = loop_back_R_0_control ? 1'h1 : _GEN_44; // @[LoopBlock.scala 903:56]
  assign _GEN_106 = loop_back_R_0_control ? 1'h1 : _GEN_46; // @[LoopBlock.scala 903:56]
  assign _GEN_107 = loop_back_R_0_control ? 1'h1 : _GEN_48; // @[LoopBlock.scala 903:56]
  assign _GEN_108 = loop_back_R_0_control ? 1'h0 : _GEN_5; // @[LoopBlock.scala 903:56]
  assign _GEN_109 = loop_back_R_0_control ? 10'h0 : _GEN_4; // @[LoopBlock.scala 903:56]
  assign _GEN_110 = loop_back_R_0_control ? 1'h0 : _GEN_6; // @[LoopBlock.scala 903:56]
  assign _GEN_111 = loop_back_R_0_control ? 1'h0 : _GEN_8; // @[LoopBlock.scala 903:56]
  assign _GEN_113 = loop_back_R_0_control ? 1'h0 : _GEN_9; // @[LoopBlock.scala 903:56]
  assign _GEN_114 = loop_back_R_0_control ? 1'h0 : _GEN_33; // @[LoopBlock.scala 903:56]
  assign _GEN_115 = loop_back_R_0_control ? 2'h1 : _GEN_89; // @[LoopBlock.scala 903:56]
  assign _GEN_116 = loop_back_R_0_control ? _GEN_36 : _GEN_82; // @[LoopBlock.scala 903:56]
  assign _GEN_117 = loop_back_R_0_control ? loop_exit_R_0_control : _GEN_87; // @[LoopBlock.scala 903:56]
  assign _GEN_118 = loop_back_R_0_control ? loop_exit_R_0_taskID : _GEN_88; // @[LoopBlock.scala 903:56]
  assign _GEN_119 = _T_662 ? _GEN_90 : active_loop_start_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_120 = _T_662 ? _GEN_91 : active_loop_start_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_121 = _T_662 ? _GEN_92 : _GEN_34; // @[LoopBlock.scala 900:55]
  assign _GEN_122 = _T_662 ? _GEN_93 : active_loop_back_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_123 = _T_662 ? _GEN_94 : active_loop_back_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_124 = _T_662 ? _GEN_95 : _GEN_35; // @[LoopBlock.scala 900:55]
  assign _GEN_125 = _T_662 ? _GEN_96 : _GEN_39; // @[LoopBlock.scala 900:55]
  assign _GEN_126 = _T_662 ? _GEN_97 : _GEN_41; // @[LoopBlock.scala 900:55]
  assign _GEN_127 = _T_662 ? _GEN_98 : _GEN_43; // @[LoopBlock.scala 900:55]
  assign _GEN_128 = _T_662 ? _GEN_99 : _GEN_45; // @[LoopBlock.scala 900:55]
  assign _GEN_129 = _T_662 ? _GEN_100 : _GEN_47; // @[LoopBlock.scala 900:55]
  assign _GEN_131 = _T_662 ? _GEN_102 : _GEN_38; // @[LoopBlock.scala 900:55]
  assign _GEN_132 = _T_662 ? _GEN_103 : _GEN_40; // @[LoopBlock.scala 900:55]
  assign _GEN_133 = _T_662 ? _GEN_104 : _GEN_42; // @[LoopBlock.scala 900:55]
  assign _GEN_134 = _T_662 ? _GEN_105 : _GEN_44; // @[LoopBlock.scala 900:55]
  assign _GEN_135 = _T_662 ? _GEN_106 : _GEN_46; // @[LoopBlock.scala 900:55]
  assign _GEN_136 = _T_662 ? _GEN_107 : _GEN_48; // @[LoopBlock.scala 900:55]
  assign _GEN_137 = _T_662 ? _GEN_108 : _GEN_5; // @[LoopBlock.scala 900:55]
  assign _GEN_138 = _T_662 ? _GEN_109 : _GEN_4; // @[LoopBlock.scala 900:55]
  assign _GEN_139 = _T_662 ? _GEN_110 : _GEN_6; // @[LoopBlock.scala 900:55]
  assign _GEN_140 = _T_662 ? _GEN_111 : _GEN_8; // @[LoopBlock.scala 900:55]
  assign _GEN_142 = _T_662 ? _GEN_113 : _GEN_9; // @[LoopBlock.scala 900:55]
  assign _GEN_143 = _T_662 ? _GEN_114 : _GEN_33; // @[LoopBlock.scala 900:55]
  assign _GEN_144 = _T_662 ? _GEN_115 : state; // @[LoopBlock.scala 900:55]
  assign _GEN_145 = _T_662 ? _GEN_116 : _GEN_36; // @[LoopBlock.scala 900:55]
  assign _GEN_146 = _T_662 ? _GEN_117 : loop_exit_R_0_control; // @[LoopBlock.scala 900:55]
  assign _GEN_147 = _T_662 ? _GEN_118 : loop_exit_R_0_taskID; // @[LoopBlock.scala 900:55]
  assign _T_711 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_148 = loop_exit_fire_R_0 ? 10'h0 : _GEN_1; // @[LoopBlock.scala 955:48]
  assign _GEN_149 = loop_exit_fire_R_0 ? 1'h0 : _GEN_2; // @[LoopBlock.scala 955:48]
  assign _GEN_150 = loop_exit_fire_R_0 ? 1'h0 : _GEN_3; // @[LoopBlock.scala 955:48]
  assign _GEN_151 = loop_exit_fire_R_0 ? 1'h0 : _GEN_5; // @[LoopBlock.scala 955:48]
  assign _GEN_152 = loop_exit_fire_R_0 ? 10'h0 : _GEN_4; // @[LoopBlock.scala 955:48]
  assign _GEN_153 = loop_exit_fire_R_0 ? 1'h0 : _GEN_6; // @[LoopBlock.scala 955:48]
  assign _GEN_154 = loop_exit_fire_R_0 ? 1'h0 : _GEN_8; // @[LoopBlock.scala 955:48]
  assign _GEN_156 = loop_exit_fire_R_0 ? 1'h0 : _GEN_9; // @[LoopBlock.scala 955:48]
  assign _GEN_157 = loop_exit_fire_R_0 ? 32'h0 : _GEN_12; // @[LoopBlock.scala 955:48]
  assign _GEN_160 = loop_exit_fire_R_0 ? 32'h0 : _GEN_16; // @[LoopBlock.scala 955:48]
  assign _GEN_161 = loop_exit_fire_R_0 ? 10'h0 : _GEN_15; // @[LoopBlock.scala 955:48]
  assign _GEN_163 = loop_exit_fire_R_0 ? 32'h0 : _GEN_20; // @[LoopBlock.scala 955:48]
  assign _GEN_164 = loop_exit_fire_R_0 ? 10'h0 : _GEN_19; // @[LoopBlock.scala 955:48]
  assign _GEN_166 = loop_exit_fire_R_0 ? 32'h0 : _GEN_24; // @[LoopBlock.scala 955:48]
  assign _GEN_167 = loop_exit_fire_R_0 ? 10'h0 : _GEN_23; // @[LoopBlock.scala 955:48]
  assign _GEN_169 = loop_exit_fire_R_0 ? 32'h0 : _GEN_28; // @[LoopBlock.scala 955:48]
  assign _GEN_172 = loop_exit_fire_R_0 ? 1'h0 : _GEN_13; // @[LoopBlock.scala 955:48]
  assign _GEN_173 = loop_exit_fire_R_0 ? 1'h0 : _GEN_17; // @[LoopBlock.scala 955:48]
  assign _GEN_174 = loop_exit_fire_R_0 ? 1'h0 : _GEN_21; // @[LoopBlock.scala 955:48]
  assign _GEN_175 = loop_exit_fire_R_0 ? 1'h0 : _GEN_25; // @[LoopBlock.scala 955:48]
  assign _GEN_176 = loop_exit_fire_R_0 ? 1'h0 : _GEN_29; // @[LoopBlock.scala 955:48]
  assign _GEN_177 = loop_exit_fire_R_0 ? 1'h0 : _GEN_33; // @[LoopBlock.scala 955:48]
  assign _GEN_178 = loop_exit_fire_R_0 ? 2'h0 : state; // @[LoopBlock.scala 955:48]
  assign _GEN_179 = _T_711 ? _GEN_148 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_180 = _T_711 ? _GEN_149 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_181 = _T_711 ? _GEN_150 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_182 = _T_711 ? _GEN_151 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_183 = _T_711 ? _GEN_152 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_184 = _T_711 ? _GEN_153 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_185 = _T_711 ? _GEN_154 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_187 = _T_711 ? _GEN_156 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_188 = _T_711 ? _GEN_157 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_191 = _T_711 ? _GEN_160 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_192 = _T_711 ? _GEN_161 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_194 = _T_711 ? _GEN_163 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_195 = _T_711 ? _GEN_164 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_197 = _T_711 ? _GEN_166 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_198 = _T_711 ? _GEN_167 : _GEN_23; // @[Conditional.scala 39:67]
  assign _GEN_200 = _T_711 ? _GEN_169 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_203 = _T_711 ? _GEN_172 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_204 = _T_711 ? _GEN_173 : _GEN_17; // @[Conditional.scala 39:67]
  assign _GEN_205 = _T_711 ? _GEN_174 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_206 = _T_711 ? _GEN_175 : _GEN_25; // @[Conditional.scala 39:67]
  assign _GEN_207 = _T_711 ? _GEN_176 : _GEN_29; // @[Conditional.scala 39:67]
  assign _GEN_208 = _T_711 ? _GEN_177 : _GEN_33; // @[Conditional.scala 39:67]
  assign _GEN_209 = _T_711 ? _GEN_178 : state; // @[Conditional.scala 39:67]
  assign _GEN_210 = _T_654 ? _GEN_119 : active_loop_start_R_control; // @[Conditional.scala 39:67]
  assign _GEN_211 = _T_654 ? _GEN_120 : active_loop_start_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_212 = _T_654 ? _GEN_121 : _GEN_34; // @[Conditional.scala 39:67]
  assign _GEN_213 = _T_654 ? _GEN_122 : active_loop_back_R_control; // @[Conditional.scala 39:67]
  assign _GEN_214 = _T_654 ? _GEN_123 : active_loop_back_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_215 = _T_654 ? _GEN_124 : _GEN_35; // @[Conditional.scala 39:67]
  assign _GEN_216 = _T_654 ? _GEN_125 : _GEN_39; // @[Conditional.scala 39:67]
  assign _GEN_217 = _T_654 ? _GEN_126 : _GEN_41; // @[Conditional.scala 39:67]
  assign _GEN_218 = _T_654 ? _GEN_127 : _GEN_43; // @[Conditional.scala 39:67]
  assign _GEN_219 = _T_654 ? _GEN_128 : _GEN_45; // @[Conditional.scala 39:67]
  assign _GEN_220 = _T_654 ? _GEN_129 : _GEN_47; // @[Conditional.scala 39:67]
  assign _GEN_222 = _T_654 ? _GEN_131 : _GEN_38; // @[Conditional.scala 39:67]
  assign _GEN_223 = _T_654 ? _GEN_132 : _GEN_40; // @[Conditional.scala 39:67]
  assign _GEN_224 = _T_654 ? _GEN_133 : _GEN_42; // @[Conditional.scala 39:67]
  assign _GEN_225 = _T_654 ? _GEN_134 : _GEN_44; // @[Conditional.scala 39:67]
  assign _GEN_226 = _T_654 ? _GEN_135 : _GEN_46; // @[Conditional.scala 39:67]
  assign _GEN_227 = _T_654 ? _GEN_136 : _GEN_48; // @[Conditional.scala 39:67]
  assign _GEN_228 = _T_654 ? _GEN_137 : _GEN_182; // @[Conditional.scala 39:67]
  assign _GEN_229 = _T_654 ? _GEN_138 : _GEN_183; // @[Conditional.scala 39:67]
  assign _GEN_230 = _T_654 ? _GEN_139 : _GEN_184; // @[Conditional.scala 39:67]
  assign _GEN_231 = _T_654 ? _GEN_140 : _GEN_185; // @[Conditional.scala 39:67]
  assign _GEN_233 = _T_654 ? _GEN_142 : _GEN_187; // @[Conditional.scala 39:67]
  assign _GEN_234 = _T_654 ? _GEN_143 : _GEN_208; // @[Conditional.scala 39:67]
  assign _GEN_235 = _T_654 ? _GEN_144 : _GEN_209; // @[Conditional.scala 39:67]
  assign _GEN_236 = _T_654 ? _GEN_145 : _GEN_36; // @[Conditional.scala 39:67]
  assign _GEN_237 = _T_654 ? _GEN_146 : loop_exit_R_0_control; // @[Conditional.scala 39:67]
  assign _GEN_238 = _T_654 ? _GEN_147 : loop_exit_R_0_taskID; // @[Conditional.scala 39:67]
  assign _GEN_239 = _T_654 ? _GEN_1 : _GEN_179; // @[Conditional.scala 39:67]
  assign _GEN_240 = _T_654 ? _GEN_2 : _GEN_180; // @[Conditional.scala 39:67]
  assign _GEN_241 = _T_654 ? _GEN_3 : _GEN_181; // @[Conditional.scala 39:67]
  assign _GEN_242 = _T_654 ? _GEN_12 : _GEN_188; // @[Conditional.scala 39:67]
  assign _GEN_245 = _T_654 ? _GEN_16 : _GEN_191; // @[Conditional.scala 39:67]
  assign _GEN_246 = _T_654 ? _GEN_15 : _GEN_192; // @[Conditional.scala 39:67]
  assign _GEN_248 = _T_654 ? _GEN_20 : _GEN_194; // @[Conditional.scala 39:67]
  assign _GEN_249 = _T_654 ? _GEN_19 : _GEN_195; // @[Conditional.scala 39:67]
  assign _GEN_251 = _T_654 ? _GEN_24 : _GEN_197; // @[Conditional.scala 39:67]
  assign _GEN_252 = _T_654 ? _GEN_23 : _GEN_198; // @[Conditional.scala 39:67]
  assign _GEN_254 = _T_654 ? _GEN_28 : _GEN_200; // @[Conditional.scala 39:67]
  assign _GEN_257 = _T_654 ? _GEN_13 : _GEN_203; // @[Conditional.scala 39:67]
  assign _GEN_258 = _T_654 ? _GEN_17 : _GEN_204; // @[Conditional.scala 39:67]
  assign _GEN_259 = _T_654 ? _GEN_21 : _GEN_205; // @[Conditional.scala 39:67]
  assign _GEN_260 = _T_654 ? _GEN_25 : _GEN_206; // @[Conditional.scala 39:67]
  assign _GEN_261 = _T_654 ? _GEN_29 : _GEN_207; // @[Conditional.scala 39:67]
  assign _GEN_262 = _T_629 ? _GEN_66 : _GEN_222; // @[Conditional.scala 40:58]
  assign _GEN_263 = _T_629 ? _GEN_67 : _GEN_223; // @[Conditional.scala 40:58]
  assign _GEN_264 = _T_629 ? _GEN_68 : _GEN_224; // @[Conditional.scala 40:58]
  assign _GEN_265 = _T_629 ? _GEN_69 : _GEN_225; // @[Conditional.scala 40:58]
  assign _GEN_266 = _T_629 ? _GEN_70 : _GEN_226; // @[Conditional.scala 40:58]
  assign _GEN_267 = _T_629 ? _GEN_71 : _GEN_227; // @[Conditional.scala 40:58]
  assign _GEN_268 = _T_629 ? _GEN_72 : _GEN_210; // @[Conditional.scala 40:58]
  assign _GEN_269 = _T_629 ? _GEN_73 : _GEN_211; // @[Conditional.scala 40:58]
  assign _GEN_270 = _T_629 ? _GEN_74 : _GEN_212; // @[Conditional.scala 40:58]
  assign _GEN_271 = _T_629 ? _GEN_75 : _GEN_213; // @[Conditional.scala 40:58]
  assign _GEN_272 = _T_629 ? _GEN_76 : _GEN_214; // @[Conditional.scala 40:58]
  assign _GEN_273 = _T_629 ? _GEN_77 : _GEN_215; // @[Conditional.scala 40:58]
  assign _GEN_274 = _T_629 ? _GEN_78 : _GEN_235; // @[Conditional.scala 40:58]
  assign _GEN_275 = _T_629 ? _GEN_79 : _GEN_237; // @[Conditional.scala 40:58]
  assign _GEN_276 = _T_629 ? _GEN_80 : _GEN_238; // @[Conditional.scala 40:58]
  assign _GEN_277 = _T_629 ? _GEN_81 : _GEN_236; // @[Conditional.scala 40:58]
  assign _GEN_278 = _T_629 ? _GEN_39 : _GEN_216; // @[Conditional.scala 40:58]
  assign _GEN_279 = _T_629 ? _GEN_41 : _GEN_217; // @[Conditional.scala 40:58]
  assign _GEN_280 = _T_629 ? _GEN_43 : _GEN_218; // @[Conditional.scala 40:58]
  assign _GEN_281 = _T_629 ? _GEN_45 : _GEN_219; // @[Conditional.scala 40:58]
  assign _GEN_282 = _T_629 ? _GEN_47 : _GEN_220; // @[Conditional.scala 40:58]
  assign _GEN_284 = _T_629 ? _GEN_5 : _GEN_228; // @[Conditional.scala 40:58]
  assign _GEN_285 = _T_629 ? _GEN_4 : _GEN_229; // @[Conditional.scala 40:58]
  assign _GEN_286 = _T_629 ? _GEN_6 : _GEN_230; // @[Conditional.scala 40:58]
  assign _GEN_287 = _T_629 ? _GEN_8 : _GEN_231; // @[Conditional.scala 40:58]
  assign _GEN_289 = _T_629 ? _GEN_9 : _GEN_233; // @[Conditional.scala 40:58]
  assign _GEN_290 = _T_629 ? _GEN_33 : _GEN_234; // @[Conditional.scala 40:58]
  assign _GEN_291 = _T_629 ? _GEN_1 : _GEN_239; // @[Conditional.scala 40:58]
  assign _GEN_292 = _T_629 ? _GEN_2 : _GEN_240; // @[Conditional.scala 40:58]
  assign _GEN_293 = _T_629 ? _GEN_3 : _GEN_241; // @[Conditional.scala 40:58]
  assign _GEN_294 = _T_629 ? _GEN_12 : _GEN_242; // @[Conditional.scala 40:58]
  assign _GEN_297 = _T_629 ? _GEN_16 : _GEN_245; // @[Conditional.scala 40:58]
  assign _GEN_298 = _T_629 ? _GEN_15 : _GEN_246; // @[Conditional.scala 40:58]
  assign _GEN_300 = _T_629 ? _GEN_20 : _GEN_248; // @[Conditional.scala 40:58]
  assign _GEN_301 = _T_629 ? _GEN_19 : _GEN_249; // @[Conditional.scala 40:58]
  assign _GEN_303 = _T_629 ? _GEN_24 : _GEN_251; // @[Conditional.scala 40:58]
  assign _GEN_304 = _T_629 ? _GEN_23 : _GEN_252; // @[Conditional.scala 40:58]
  assign _GEN_306 = _T_629 ? _GEN_28 : _GEN_254; // @[Conditional.scala 40:58]
  assign _GEN_309 = _T_629 ? _GEN_13 : _GEN_257; // @[Conditional.scala 40:58]
  assign _GEN_310 = _T_629 ? _GEN_17 : _GEN_258; // @[Conditional.scala 40:58]
  assign _GEN_311 = _T_629 ? _GEN_21 : _GEN_259; // @[Conditional.scala 40:58]
  assign _GEN_312 = _T_629 ? _GEN_25 : _GEN_260; // @[Conditional.scala 40:58]
  assign _GEN_313 = _T_629 ? _GEN_29 : _GEN_261; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_taskID = in_live_in_R_3_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_taskID = _RAND_13[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_21[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_35[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_38[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_41[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  state = _RAND_45[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_577) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_654) begin
          if (_T_577) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_577) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_577) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_577) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_654) begin
          if (_T_577) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_577) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_577) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_577) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_577) begin
            enable_valid_R <= 1'h1;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_577) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_577) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_580) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_580) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_580) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_580) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_580) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_580) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_580) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_580) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_580) begin
          loop_back_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_580) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_580) begin
              loop_back_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_580) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_583) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_583) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_583) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_583) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_8;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_583) begin
          loop_finish_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_583) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_583) begin
              loop_finish_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_583) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_629) begin
        if (_T_586) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_654) begin
          if (_T_586) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_586) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_586) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_589) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_654) begin
          if (_T_589) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_taskID <= 10'h0;
            end else begin
              if (_T_589) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_589) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_629) begin
        if (_T_589) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_654) begin
          if (_T_589) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_589) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_589) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_592) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_654) begin
          if (_T_592) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_taskID <= 10'h0;
            end else begin
              if (_T_592) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_592) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_629) begin
        if (_T_592) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_654) begin
          if (_T_592) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_592) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_592) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_595) begin
          in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
        end
      end else begin
        if (_T_654) begin
          if (_T_595) begin
            in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_taskID <= 10'h0;
            end else begin
              if (_T_595) begin
                in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
              end
            end
          end else begin
            if (_T_595) begin
              in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_629) begin
        if (_T_595) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_654) begin
          if (_T_595) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_595) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_595) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_629) begin
        if (_T_598) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_654) begin
          if (_T_598) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_598) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_598) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_586) begin
          in_live_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_586) begin
            in_live_in_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_586) begin
                in_live_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_586) begin
              in_live_in_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_589) begin
          in_live_in_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_589) begin
            in_live_in_valid_R_1 <= 1'h1;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              if (_T_589) begin
                in_live_in_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_589) begin
              in_live_in_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_592) begin
          in_live_in_valid_R_2 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_592) begin
            in_live_in_valid_R_2 <= 1'h1;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              if (_T_592) begin
                in_live_in_valid_R_2 <= 1'h1;
              end
            end
          end else begin
            if (_T_592) begin
              in_live_in_valid_R_2 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_595) begin
          in_live_in_valid_R_3 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_595) begin
            in_live_in_valid_R_3 <= 1'h1;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              if (_T_595) begin
                in_live_in_valid_R_3 <= 1'h1;
              end
            end
          end else begin
            if (_T_595) begin
              in_live_in_valid_R_3 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_598) begin
          in_live_in_valid_R_4 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_598) begin
            in_live_in_valid_R_4 <= 1'h1;
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              if (_T_598) begin
                in_live_in_valid_R_4 <= 1'h1;
              end
            end
          end else begin
            if (_T_598) begin
              in_live_in_valid_R_4 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_601) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_601) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_601) begin
          in_carry_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_601) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_601) begin
              in_carry_in_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_601) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            out_live_in_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_610) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_610) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_610) begin
                out_live_in_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_610) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_0_0 <= _GEN_38;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            out_live_in_valid_R_1_0 <= 1'h1;
          end else begin
            if (_T_613) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_613) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_1_0 <= 1'h1;
            end else begin
              if (_T_613) begin
                out_live_in_valid_R_1_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_613) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_1_0 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            out_live_in_valid_R_2_0 <= 1'h1;
          end else begin
            if (_T_616) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_616) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_2_0 <= 1'h1;
            end else begin
              if (_T_616) begin
                out_live_in_valid_R_2_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_616) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_2_0 <= _GEN_42;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            out_live_in_valid_R_3_0 <= 1'h1;
          end else begin
            if (_T_619) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_619) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_3_0 <= 1'h1;
            end else begin
              if (_T_619) begin
                out_live_in_valid_R_3_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_619) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_3_0 <= _GEN_44;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            out_live_in_valid_R_4_0 <= 1'h1;
          end else begin
            if (_T_622) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_622) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_4_0 <= 1'h1;
            end else begin
              if (_T_622) begin
                out_live_in_valid_R_4_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_622) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_4_0 <= _GEN_46;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_610) begin
          out_live_in_fire_R_0_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              if (_T_610) begin
                out_live_in_fire_R_0_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_610) begin
              out_live_in_fire_R_0_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_610) begin
            out_live_in_fire_R_0_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_613) begin
          out_live_in_fire_R_1_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              if (_T_613) begin
                out_live_in_fire_R_1_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_613) begin
              out_live_in_fire_R_1_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_613) begin
            out_live_in_fire_R_1_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_616) begin
          out_live_in_fire_R_2_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              if (_T_616) begin
                out_live_in_fire_R_2_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_616) begin
              out_live_in_fire_R_2_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_616) begin
            out_live_in_fire_R_2_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_619) begin
          out_live_in_fire_R_3_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              if (_T_619) begin
                out_live_in_fire_R_3_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_619) begin
              out_live_in_fire_R_3_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_619) begin
            out_live_in_fire_R_3_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_622) begin
          out_live_in_fire_R_4_0 <= 1'h1;
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              if (_T_622) begin
                out_live_in_fire_R_4_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_622) begin
              out_live_in_fire_R_4_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_622) begin
            out_live_in_fire_R_4_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            out_carry_out_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_625) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_625) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              out_carry_out_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_625) begin
                out_carry_out_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_625) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_carry_out_valid_R_0_0 <= _GEN_48;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            active_loop_start_R_control <= 1'h1;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            active_loop_start_valid_R <= 1'h1;
          end else begin
            if (_T_603) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_603) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              active_loop_start_valid_R <= 1'h1;
            end else begin
              if (_T_603) begin
                active_loop_start_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_603) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_start_valid_R <= _GEN_34;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_control <= 1'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            active_loop_back_valid_R <= 1'h1;
          end else begin
            if (_T_605) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_605) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              active_loop_back_valid_R <= 1'h1;
            end else begin
              if (_T_605) begin
                active_loop_back_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_605) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_back_valid_R <= _GEN_35;
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 10'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 10'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_control <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_control <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            if (_T_607) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_607) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              if (_T_607) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              if (loop_finish_R_0_control) begin
                loop_exit_valid_R_0 <= 1'h1;
              end else begin
                if (_T_607) begin
                  loop_exit_valid_R_0 <= 1'h0;
                end
              end
            end
          end else begin
            loop_exit_valid_R_0 <= _GEN_36;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_36;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      if (_T_607) begin
        loop_exit_fire_R_0 <= 1'h1;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_629) begin
        if (_T_634) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_654) begin
          if (_T_662) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_711) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [9:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [9:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [9:0]  io_InLiveIn_3_bits_taskID,
  input  [31:0] io_InLiveIn_3_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [9:0]  io_OutLiveIn_field3_0_bits_taskID,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [9:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [9:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [9:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [9:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [9:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [9:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [9:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [9:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_2;
  reg [9:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_3;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_5;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_6;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_7;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_8;
  reg [9:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [9:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [9:0] in_live_in_R_3_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_15;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_16;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_17;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_18;
  reg [9:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_19;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_20;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_21;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_22;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_23;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_24;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_25;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_26;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_29;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_30;
  reg [9:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_31;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_32;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_33;
  reg [9:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_34;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_35;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_36;
  reg [9:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_37;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_38;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_39;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_40;
  wire  _T_519; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[LoopBlock.scala 596:26]
  wire  _GEN_2; // @[LoopBlock.scala 596:26]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_522; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_4; // @[LoopBlock.scala 603:33]
  wire  _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_525; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_528; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[LoopBlock.scala 623:33]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_531; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_15; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_16; // @[LoopBlock.scala 623:33]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_534; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_19; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_20; // @[LoopBlock.scala 623:33]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_537; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_23; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_24; // @[LoopBlock.scala 623:33]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_540; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_27; // @[LoopBlock.scala 641:37]
  wire [31:0] _GEN_28; // @[LoopBlock.scala 641:37]
  wire  _GEN_29; // @[LoopBlock.scala 641:37]
  wire  _T_542; // @[Decoupled.scala 37:37]
  wire  _GEN_30; // @[LoopBlock.scala 704:39]
  wire  _T_544; // @[Decoupled.scala 37:37]
  wire  _GEN_31; // @[LoopBlock.scala 708:38]
  wire  _T_546; // @[Decoupled.scala 37:37]
  wire  _GEN_32; // @[LoopBlock.scala 713:33]
  wire  _GEN_33; // @[LoopBlock.scala 713:33]
  wire  _T_549; // @[Decoupled.scala 37:37]
  wire  _GEN_34; // @[LoopBlock.scala 722:57]
  wire  _GEN_35; // @[LoopBlock.scala 722:57]
  wire  _T_552; // @[Decoupled.scala 37:37]
  wire  _GEN_36; // @[LoopBlock.scala 722:57]
  wire  _GEN_37; // @[LoopBlock.scala 722:57]
  wire  _T_555; // @[Decoupled.scala 37:37]
  wire  _GEN_38; // @[LoopBlock.scala 722:57]
  wire  _GEN_39; // @[LoopBlock.scala 722:57]
  wire  _T_558; // @[Decoupled.scala 37:37]
  wire  _GEN_40; // @[LoopBlock.scala 722:57]
  wire  _GEN_41; // @[LoopBlock.scala 722:57]
  wire  _T_561; // @[Decoupled.scala 37:37]
  wire  _GEN_42; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_41;
  wire  _T_565; // @[Conditional.scala 37:30]
  wire  _T_566; // @[LoopBlock.scala 765:35]
  wire  _T_567; // @[LoopBlock.scala 765:35]
  wire  _T_568; // @[LoopBlock.scala 765:35]
  wire  _T_569; // @[LoopBlock.scala 869:28]
  wire  _GEN_44; // @[LoopBlock.scala 870:26]
  wire  _GEN_45; // @[LoopBlock.scala 870:26]
  wire  _GEN_46; // @[LoopBlock.scala 870:26]
  wire  _GEN_47; // @[LoopBlock.scala 870:26]
  wire  _GEN_48; // @[LoopBlock.scala 870:26]
  wire  _GEN_49; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_50; // @[LoopBlock.scala 870:26]
  wire  _GEN_51; // @[LoopBlock.scala 870:26]
  wire  _GEN_52; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_53; // @[LoopBlock.scala 870:26]
  wire  _GEN_54; // @[LoopBlock.scala 870:26]
  wire [1:0] _GEN_55; // @[LoopBlock.scala 870:26]
  wire  _GEN_56; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_57; // @[LoopBlock.scala 870:26]
  wire  _GEN_58; // @[LoopBlock.scala 870:26]
  wire  _GEN_59; // @[LoopBlock.scala 869:48]
  wire  _GEN_60; // @[LoopBlock.scala 869:48]
  wire  _GEN_61; // @[LoopBlock.scala 869:48]
  wire  _GEN_62; // @[LoopBlock.scala 869:48]
  wire  _GEN_63; // @[LoopBlock.scala 869:48]
  wire  _GEN_64; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_65; // @[LoopBlock.scala 869:48]
  wire  _GEN_66; // @[LoopBlock.scala 869:48]
  wire  _GEN_67; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_68; // @[LoopBlock.scala 869:48]
  wire  _GEN_69; // @[LoopBlock.scala 869:48]
  wire [1:0] _GEN_70; // @[LoopBlock.scala 869:48]
  wire  _GEN_71; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_72; // @[LoopBlock.scala 869:48]
  wire  _GEN_73; // @[LoopBlock.scala 869:48]
  wire  _T_588; // @[Conditional.scala 37:30]
  wire  _T_589; // @[LoopBlock.scala 898:30]
  wire  _T_592; // @[LoopBlock.scala 828:26]
  wire  _T_593; // @[LoopBlock.scala 828:26]
  wire  _T_594; // @[LoopBlock.scala 828:26]
  wire  _T_595; // @[LoopBlock.scala 899:29]
  wire  _GEN_74; // @[LoopBlock.scala 936:64]
  wire  _GEN_75; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_76; // @[LoopBlock.scala 936:64]
  wire  _GEN_77; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_78; // @[LoopBlock.scala 936:64]
  wire  _GEN_79; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_80; // @[LoopBlock.scala 936:64]
  wire [1:0] _GEN_81; // @[LoopBlock.scala 936:64]
  wire  _GEN_82; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_83; // @[LoopBlock.scala 903:56]
  wire  _GEN_84; // @[LoopBlock.scala 903:56]
  wire  _GEN_85; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_86; // @[LoopBlock.scala 903:56]
  wire  _GEN_87; // @[LoopBlock.scala 903:56]
  wire  _GEN_88; // @[LoopBlock.scala 903:56]
  wire  _GEN_89; // @[LoopBlock.scala 903:56]
  wire  _GEN_90; // @[LoopBlock.scala 903:56]
  wire  _GEN_91; // @[LoopBlock.scala 903:56]
  wire  _GEN_93; // @[LoopBlock.scala 903:56]
  wire  _GEN_94; // @[LoopBlock.scala 903:56]
  wire  _GEN_95; // @[LoopBlock.scala 903:56]
  wire  _GEN_96; // @[LoopBlock.scala 903:56]
  wire  _GEN_97; // @[LoopBlock.scala 903:56]
  wire  _GEN_98; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_99; // @[LoopBlock.scala 903:56]
  wire  _GEN_100; // @[LoopBlock.scala 903:56]
  wire  _GEN_101; // @[LoopBlock.scala 903:56]
  wire  _GEN_103; // @[LoopBlock.scala 903:56]
  wire  _GEN_104; // @[LoopBlock.scala 903:56]
  wire [1:0] _GEN_105; // @[LoopBlock.scala 903:56]
  wire  _GEN_106; // @[LoopBlock.scala 903:56]
  wire  _GEN_107; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_108; // @[LoopBlock.scala 903:56]
  wire  _GEN_109; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_110; // @[LoopBlock.scala 900:55]
  wire  _GEN_111; // @[LoopBlock.scala 900:55]
  wire  _GEN_112; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_113; // @[LoopBlock.scala 900:55]
  wire  _GEN_114; // @[LoopBlock.scala 900:55]
  wire  _GEN_115; // @[LoopBlock.scala 900:55]
  wire  _GEN_116; // @[LoopBlock.scala 900:55]
  wire  _GEN_117; // @[LoopBlock.scala 900:55]
  wire  _GEN_118; // @[LoopBlock.scala 900:55]
  wire  _GEN_120; // @[LoopBlock.scala 900:55]
  wire  _GEN_121; // @[LoopBlock.scala 900:55]
  wire  _GEN_122; // @[LoopBlock.scala 900:55]
  wire  _GEN_123; // @[LoopBlock.scala 900:55]
  wire  _GEN_124; // @[LoopBlock.scala 900:55]
  wire  _GEN_125; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_126; // @[LoopBlock.scala 900:55]
  wire  _GEN_127; // @[LoopBlock.scala 900:55]
  wire  _GEN_128; // @[LoopBlock.scala 900:55]
  wire  _GEN_130; // @[LoopBlock.scala 900:55]
  wire  _GEN_131; // @[LoopBlock.scala 900:55]
  wire [1:0] _GEN_132; // @[LoopBlock.scala 900:55]
  wire  _GEN_133; // @[LoopBlock.scala 900:55]
  wire  _GEN_134; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_135; // @[LoopBlock.scala 900:55]
  wire  _T_642; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_136; // @[LoopBlock.scala 955:48]
  wire  _GEN_137; // @[LoopBlock.scala 955:48]
  wire  _GEN_138; // @[LoopBlock.scala 955:48]
  wire  _GEN_139; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_140; // @[LoopBlock.scala 955:48]
  wire  _GEN_141; // @[LoopBlock.scala 955:48]
  wire  _GEN_142; // @[LoopBlock.scala 955:48]
  wire  _GEN_144; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_145; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_148; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_149; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_151; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_152; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_154; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_155; // @[LoopBlock.scala 955:48]
  wire  _GEN_157; // @[LoopBlock.scala 955:48]
  wire  _GEN_158; // @[LoopBlock.scala 955:48]
  wire  _GEN_159; // @[LoopBlock.scala 955:48]
  wire  _GEN_160; // @[LoopBlock.scala 955:48]
  wire  _GEN_161; // @[LoopBlock.scala 955:48]
  wire [1:0] _GEN_162; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_163; // @[Conditional.scala 39:67]
  wire  _GEN_164; // @[Conditional.scala 39:67]
  wire  _GEN_165; // @[Conditional.scala 39:67]
  wire  _GEN_166; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_167; // @[Conditional.scala 39:67]
  wire  _GEN_168; // @[Conditional.scala 39:67]
  wire  _GEN_169; // @[Conditional.scala 39:67]
  wire  _GEN_171; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_172; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_175; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_176; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_178; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_179; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_181; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_182; // @[Conditional.scala 39:67]
  wire  _GEN_184; // @[Conditional.scala 39:67]
  wire  _GEN_185; // @[Conditional.scala 39:67]
  wire  _GEN_186; // @[Conditional.scala 39:67]
  wire  _GEN_187; // @[Conditional.scala 39:67]
  wire  _GEN_188; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_189; // @[Conditional.scala 39:67]
  wire  _GEN_190; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_191; // @[Conditional.scala 39:67]
  wire  _GEN_192; // @[Conditional.scala 39:67]
  wire  _GEN_193; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_194; // @[Conditional.scala 39:67]
  wire  _GEN_195; // @[Conditional.scala 39:67]
  wire  _GEN_196; // @[Conditional.scala 39:67]
  wire  _GEN_197; // @[Conditional.scala 39:67]
  wire  _GEN_198; // @[Conditional.scala 39:67]
  wire  _GEN_199; // @[Conditional.scala 39:67]
  wire  _GEN_201; // @[Conditional.scala 39:67]
  wire  _GEN_202; // @[Conditional.scala 39:67]
  wire  _GEN_203; // @[Conditional.scala 39:67]
  wire  _GEN_204; // @[Conditional.scala 39:67]
  wire  _GEN_205; // @[Conditional.scala 39:67]
  wire  _GEN_206; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_207; // @[Conditional.scala 39:67]
  wire  _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_209; // @[Conditional.scala 39:67]
  wire  _GEN_211; // @[Conditional.scala 39:67]
  wire  _GEN_212; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_213; // @[Conditional.scala 39:67]
  wire  _GEN_214; // @[Conditional.scala 39:67]
  wire  _GEN_215; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_216; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_217; // @[Conditional.scala 39:67]
  wire  _GEN_218; // @[Conditional.scala 39:67]
  wire  _GEN_219; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_220; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_223; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_224; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_226; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_227; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_229; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_230; // @[Conditional.scala 39:67]
  wire  _GEN_232; // @[Conditional.scala 39:67]
  wire  _GEN_233; // @[Conditional.scala 39:67]
  wire  _GEN_234; // @[Conditional.scala 39:67]
  wire  _GEN_235; // @[Conditional.scala 39:67]
  wire  _GEN_236; // @[Conditional.scala 40:58]
  wire  _GEN_237; // @[Conditional.scala 40:58]
  wire  _GEN_238; // @[Conditional.scala 40:58]
  wire  _GEN_239; // @[Conditional.scala 40:58]
  wire  _GEN_240; // @[Conditional.scala 40:58]
  wire  _GEN_241; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_242; // @[Conditional.scala 40:58]
  wire  _GEN_243; // @[Conditional.scala 40:58]
  wire  _GEN_244; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_245; // @[Conditional.scala 40:58]
  wire  _GEN_246; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_247; // @[Conditional.scala 40:58]
  wire  _GEN_248; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_249; // @[Conditional.scala 40:58]
  wire  _GEN_250; // @[Conditional.scala 40:58]
  wire  _GEN_251; // @[Conditional.scala 40:58]
  wire  _GEN_252; // @[Conditional.scala 40:58]
  wire  _GEN_253; // @[Conditional.scala 40:58]
  wire  _GEN_254; // @[Conditional.scala 40:58]
  wire  _GEN_256; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_257; // @[Conditional.scala 40:58]
  wire  _GEN_258; // @[Conditional.scala 40:58]
  wire  _GEN_259; // @[Conditional.scala 40:58]
  wire  _GEN_261; // @[Conditional.scala 40:58]
  wire  _GEN_262; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_263; // @[Conditional.scala 40:58]
  wire  _GEN_264; // @[Conditional.scala 40:58]
  wire  _GEN_265; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_266; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_269; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_270; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_272; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_273; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_275; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_276; // @[Conditional.scala 40:58]
  wire  _GEN_278; // @[Conditional.scala 40:58]
  wire  _GEN_279; // @[Conditional.scala 40:58]
  wire  _GEN_280; // @[Conditional.scala 40:58]
  wire  _GEN_281; // @[Conditional.scala 40:58]
  assign _T_519 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_519 ? io_enable_bits_taskID : enable_R_taskID; // @[LoopBlock.scala 596:26]
  assign _GEN_2 = _T_519 ? io_enable_bits_control : enable_R_control; // @[LoopBlock.scala 596:26]
  assign _GEN_3 = _T_519 ? 1'h1 : enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_522 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_522 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_522 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_522 ? 1'h1 : loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_525 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_525 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_525 ? 1'h1 : loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_528 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_528 ? io_InLiveIn_0_bits_data : in_live_in_R_0_data; // @[LoopBlock.scala 623:33]
  assign _GEN_13 = _T_528 ? 1'h1 : in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_531 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_15 = _T_531 ? io_InLiveIn_1_bits_taskID : in_live_in_R_1_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_16 = _T_531 ? io_InLiveIn_1_bits_data : in_live_in_R_1_data; // @[LoopBlock.scala 623:33]
  assign _GEN_17 = _T_531 ? 1'h1 : in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_534 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_19 = _T_534 ? io_InLiveIn_2_bits_taskID : in_live_in_R_2_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_20 = _T_534 ? io_InLiveIn_2_bits_data : in_live_in_R_2_data; // @[LoopBlock.scala 623:33]
  assign _GEN_21 = _T_534 ? 1'h1 : in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_537 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_23 = _T_537 ? io_InLiveIn_3_bits_taskID : in_live_in_R_3_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_24 = _T_537 ? io_InLiveIn_3_bits_data : in_live_in_R_3_data; // @[LoopBlock.scala 623:33]
  assign _GEN_25 = _T_537 ? 1'h1 : in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_540 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_27 = _T_540 ? io_CarryDepenIn_0_bits_taskID : in_carry_in_R_0_taskID; // @[LoopBlock.scala 641:37]
  assign _GEN_28 = _T_540 ? io_CarryDepenIn_0_bits_data : in_carry_in_R_0_data; // @[LoopBlock.scala 641:37]
  assign _GEN_29 = _T_540 ? 1'h1 : in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_542 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 37:37]
  assign _GEN_30 = _T_542 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_544 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 37:37]
  assign _GEN_31 = _T_544 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_546 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_32 = _T_546 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_33 = _T_546 ? 1'h1 : loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_549 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_34 = _T_549 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_35 = _T_549 ? 1'h1 : out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_552 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_36 = _T_552 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_37 = _T_552 ? 1'h1 : out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_555 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_38 = _T_555 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_39 = _T_555 ? 1'h1 : out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_558 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_40 = _T_558 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_41 = _T_558 ? 1'h1 : out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_561 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_42 = _T_561 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_565 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_566 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_567 = _T_566 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_568 = _T_567 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_569 = _T_568 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_44 = enable_R_control ? 1'h1 : _GEN_34; // @[LoopBlock.scala 870:26]
  assign _GEN_45 = enable_R_control ? 1'h1 : _GEN_36; // @[LoopBlock.scala 870:26]
  assign _GEN_46 = enable_R_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_47 = enable_R_control ? 1'h1 : _GEN_40; // @[LoopBlock.scala 870:26]
  assign _GEN_48 = enable_R_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_49 = enable_R_control ? 1'h1 : active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_50 = enable_R_control ? enable_R_taskID : active_loop_start_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_51 = enable_R_control ? 1'h1 : _GEN_30; // @[LoopBlock.scala 870:26]
  assign _GEN_52 = enable_R_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_53 = enable_R_control ? enable_R_taskID : active_loop_back_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_54 = enable_R_control ? 1'h1 : _GEN_31; // @[LoopBlock.scala 870:26]
  assign _GEN_55 = enable_R_control ? 2'h1 : 2'h2; // @[LoopBlock.scala 870:26]
  assign _GEN_56 = enable_R_control ? loop_exit_R_0_control : 1'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_57 = enable_R_control ? loop_exit_R_0_taskID : 10'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_58 = enable_R_control ? _GEN_32 : 1'h1; // @[LoopBlock.scala 870:26]
  assign _GEN_59 = _T_569 ? _GEN_44 : _GEN_34; // @[LoopBlock.scala 869:48]
  assign _GEN_60 = _T_569 ? _GEN_45 : _GEN_36; // @[LoopBlock.scala 869:48]
  assign _GEN_61 = _T_569 ? _GEN_46 : _GEN_38; // @[LoopBlock.scala 869:48]
  assign _GEN_62 = _T_569 ? _GEN_47 : _GEN_40; // @[LoopBlock.scala 869:48]
  assign _GEN_63 = _T_569 ? _GEN_48 : _GEN_42; // @[LoopBlock.scala 869:48]
  assign _GEN_64 = _T_569 ? _GEN_49 : active_loop_start_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_65 = _T_569 ? _GEN_50 : active_loop_start_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_66 = _T_569 ? _GEN_51 : _GEN_30; // @[LoopBlock.scala 869:48]
  assign _GEN_67 = _T_569 ? _GEN_52 : active_loop_back_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_68 = _T_569 ? _GEN_53 : active_loop_back_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_69 = _T_569 ? _GEN_54 : _GEN_31; // @[LoopBlock.scala 869:48]
  assign _GEN_70 = _T_569 ? _GEN_55 : state; // @[LoopBlock.scala 869:48]
  assign _GEN_71 = _T_569 ? _GEN_56 : loop_exit_R_0_control; // @[LoopBlock.scala 869:48]
  assign _GEN_72 = _T_569 ? _GEN_57 : loop_exit_R_0_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_73 = _T_569 ? _GEN_58 : _GEN_32; // @[LoopBlock.scala 869:48]
  assign _T_588 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_589 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_592 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_593 = _T_592 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_594 = _T_593 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_595 = _T_589 & _T_594; // @[LoopBlock.scala 899:29]
  assign _GEN_74 = loop_finish_R_0_control ? 1'h1 : _GEN_32; // @[LoopBlock.scala 936:64]
  assign _GEN_75 = loop_finish_R_0_control ? 1'h0 : active_loop_start_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_76 = loop_finish_R_0_control ? 10'h0 : active_loop_start_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_77 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_78 = loop_finish_R_0_control ? 10'h0 : active_loop_back_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_79 = loop_finish_R_0_control ? 1'h1 : loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_80 = loop_finish_R_0_control ? loop_back_R_0_taskID : loop_exit_R_0_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_81 = loop_finish_R_0_control ? 2'h2 : state; // @[LoopBlock.scala 936:64]
  assign _GEN_82 = loop_back_R_0_control ? 1'h0 : _GEN_75; // @[LoopBlock.scala 903:56]
  assign _GEN_83 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_76; // @[LoopBlock.scala 903:56]
  assign _GEN_84 = loop_back_R_0_control ? 1'h1 : _GEN_30; // @[LoopBlock.scala 903:56]
  assign _GEN_85 = loop_back_R_0_control ? 1'h1 : _GEN_77; // @[LoopBlock.scala 903:56]
  assign _GEN_86 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_78; // @[LoopBlock.scala 903:56]
  assign _GEN_87 = loop_back_R_0_control ? 1'h1 : _GEN_31; // @[LoopBlock.scala 903:56]
  assign _GEN_88 = loop_back_R_0_control ? 1'h0 : _GEN_35; // @[LoopBlock.scala 903:56]
  assign _GEN_89 = loop_back_R_0_control ? 1'h0 : _GEN_37; // @[LoopBlock.scala 903:56]
  assign _GEN_90 = loop_back_R_0_control ? 1'h0 : _GEN_39; // @[LoopBlock.scala 903:56]
  assign _GEN_91 = loop_back_R_0_control ? 1'h0 : _GEN_41; // @[LoopBlock.scala 903:56]
  assign _GEN_93 = loop_back_R_0_control ? 1'h1 : _GEN_34; // @[LoopBlock.scala 903:56]
  assign _GEN_94 = loop_back_R_0_control ? 1'h1 : _GEN_36; // @[LoopBlock.scala 903:56]
  assign _GEN_95 = loop_back_R_0_control ? 1'h1 : _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_96 = loop_back_R_0_control ? 1'h1 : _GEN_40; // @[LoopBlock.scala 903:56]
  assign _GEN_97 = loop_back_R_0_control ? 1'h1 : _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_98 = loop_back_R_0_control ? 1'h0 : _GEN_5; // @[LoopBlock.scala 903:56]
  assign _GEN_99 = loop_back_R_0_control ? 10'h0 : _GEN_4; // @[LoopBlock.scala 903:56]
  assign _GEN_100 = loop_back_R_0_control ? 1'h0 : _GEN_6; // @[LoopBlock.scala 903:56]
  assign _GEN_101 = loop_back_R_0_control ? 1'h0 : _GEN_8; // @[LoopBlock.scala 903:56]
  assign _GEN_103 = loop_back_R_0_control ? 1'h0 : _GEN_9; // @[LoopBlock.scala 903:56]
  assign _GEN_104 = loop_back_R_0_control ? 1'h0 : _GEN_29; // @[LoopBlock.scala 903:56]
  assign _GEN_105 = loop_back_R_0_control ? 2'h1 : _GEN_81; // @[LoopBlock.scala 903:56]
  assign _GEN_106 = loop_back_R_0_control ? _GEN_32 : _GEN_74; // @[LoopBlock.scala 903:56]
  assign _GEN_107 = loop_back_R_0_control ? loop_exit_R_0_control : _GEN_79; // @[LoopBlock.scala 903:56]
  assign _GEN_108 = loop_back_R_0_control ? loop_exit_R_0_taskID : _GEN_80; // @[LoopBlock.scala 903:56]
  assign _GEN_109 = _T_595 ? _GEN_82 : active_loop_start_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_110 = _T_595 ? _GEN_83 : active_loop_start_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_111 = _T_595 ? _GEN_84 : _GEN_30; // @[LoopBlock.scala 900:55]
  assign _GEN_112 = _T_595 ? _GEN_85 : active_loop_back_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_113 = _T_595 ? _GEN_86 : active_loop_back_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_114 = _T_595 ? _GEN_87 : _GEN_31; // @[LoopBlock.scala 900:55]
  assign _GEN_115 = _T_595 ? _GEN_88 : _GEN_35; // @[LoopBlock.scala 900:55]
  assign _GEN_116 = _T_595 ? _GEN_89 : _GEN_37; // @[LoopBlock.scala 900:55]
  assign _GEN_117 = _T_595 ? _GEN_90 : _GEN_39; // @[LoopBlock.scala 900:55]
  assign _GEN_118 = _T_595 ? _GEN_91 : _GEN_41; // @[LoopBlock.scala 900:55]
  assign _GEN_120 = _T_595 ? _GEN_93 : _GEN_34; // @[LoopBlock.scala 900:55]
  assign _GEN_121 = _T_595 ? _GEN_94 : _GEN_36; // @[LoopBlock.scala 900:55]
  assign _GEN_122 = _T_595 ? _GEN_95 : _GEN_38; // @[LoopBlock.scala 900:55]
  assign _GEN_123 = _T_595 ? _GEN_96 : _GEN_40; // @[LoopBlock.scala 900:55]
  assign _GEN_124 = _T_595 ? _GEN_97 : _GEN_42; // @[LoopBlock.scala 900:55]
  assign _GEN_125 = _T_595 ? _GEN_98 : _GEN_5; // @[LoopBlock.scala 900:55]
  assign _GEN_126 = _T_595 ? _GEN_99 : _GEN_4; // @[LoopBlock.scala 900:55]
  assign _GEN_127 = _T_595 ? _GEN_100 : _GEN_6; // @[LoopBlock.scala 900:55]
  assign _GEN_128 = _T_595 ? _GEN_101 : _GEN_8; // @[LoopBlock.scala 900:55]
  assign _GEN_130 = _T_595 ? _GEN_103 : _GEN_9; // @[LoopBlock.scala 900:55]
  assign _GEN_131 = _T_595 ? _GEN_104 : _GEN_29; // @[LoopBlock.scala 900:55]
  assign _GEN_132 = _T_595 ? _GEN_105 : state; // @[LoopBlock.scala 900:55]
  assign _GEN_133 = _T_595 ? _GEN_106 : _GEN_32; // @[LoopBlock.scala 900:55]
  assign _GEN_134 = _T_595 ? _GEN_107 : loop_exit_R_0_control; // @[LoopBlock.scala 900:55]
  assign _GEN_135 = _T_595 ? _GEN_108 : loop_exit_R_0_taskID; // @[LoopBlock.scala 900:55]
  assign _T_642 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_136 = loop_exit_fire_R_0 ? 10'h0 : _GEN_1; // @[LoopBlock.scala 955:48]
  assign _GEN_137 = loop_exit_fire_R_0 ? 1'h0 : _GEN_2; // @[LoopBlock.scala 955:48]
  assign _GEN_138 = loop_exit_fire_R_0 ? 1'h0 : _GEN_3; // @[LoopBlock.scala 955:48]
  assign _GEN_139 = loop_exit_fire_R_0 ? 1'h0 : _GEN_5; // @[LoopBlock.scala 955:48]
  assign _GEN_140 = loop_exit_fire_R_0 ? 10'h0 : _GEN_4; // @[LoopBlock.scala 955:48]
  assign _GEN_141 = loop_exit_fire_R_0 ? 1'h0 : _GEN_6; // @[LoopBlock.scala 955:48]
  assign _GEN_142 = loop_exit_fire_R_0 ? 1'h0 : _GEN_8; // @[LoopBlock.scala 955:48]
  assign _GEN_144 = loop_exit_fire_R_0 ? 1'h0 : _GEN_9; // @[LoopBlock.scala 955:48]
  assign _GEN_145 = loop_exit_fire_R_0 ? 32'h0 : _GEN_12; // @[LoopBlock.scala 955:48]
  assign _GEN_148 = loop_exit_fire_R_0 ? 32'h0 : _GEN_16; // @[LoopBlock.scala 955:48]
  assign _GEN_149 = loop_exit_fire_R_0 ? 10'h0 : _GEN_15; // @[LoopBlock.scala 955:48]
  assign _GEN_151 = loop_exit_fire_R_0 ? 32'h0 : _GEN_20; // @[LoopBlock.scala 955:48]
  assign _GEN_152 = loop_exit_fire_R_0 ? 10'h0 : _GEN_19; // @[LoopBlock.scala 955:48]
  assign _GEN_154 = loop_exit_fire_R_0 ? 32'h0 : _GEN_24; // @[LoopBlock.scala 955:48]
  assign _GEN_155 = loop_exit_fire_R_0 ? 10'h0 : _GEN_23; // @[LoopBlock.scala 955:48]
  assign _GEN_157 = loop_exit_fire_R_0 ? 1'h0 : _GEN_13; // @[LoopBlock.scala 955:48]
  assign _GEN_158 = loop_exit_fire_R_0 ? 1'h0 : _GEN_17; // @[LoopBlock.scala 955:48]
  assign _GEN_159 = loop_exit_fire_R_0 ? 1'h0 : _GEN_21; // @[LoopBlock.scala 955:48]
  assign _GEN_160 = loop_exit_fire_R_0 ? 1'h0 : _GEN_25; // @[LoopBlock.scala 955:48]
  assign _GEN_161 = loop_exit_fire_R_0 ? 1'h0 : _GEN_29; // @[LoopBlock.scala 955:48]
  assign _GEN_162 = loop_exit_fire_R_0 ? 2'h0 : state; // @[LoopBlock.scala 955:48]
  assign _GEN_163 = _T_642 ? _GEN_136 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_164 = _T_642 ? _GEN_137 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_165 = _T_642 ? _GEN_138 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_166 = _T_642 ? _GEN_139 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_167 = _T_642 ? _GEN_140 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_168 = _T_642 ? _GEN_141 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_169 = _T_642 ? _GEN_142 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_171 = _T_642 ? _GEN_144 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_172 = _T_642 ? _GEN_145 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_175 = _T_642 ? _GEN_148 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_176 = _T_642 ? _GEN_149 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_178 = _T_642 ? _GEN_151 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_179 = _T_642 ? _GEN_152 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_181 = _T_642 ? _GEN_154 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_182 = _T_642 ? _GEN_155 : _GEN_23; // @[Conditional.scala 39:67]
  assign _GEN_184 = _T_642 ? _GEN_157 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_185 = _T_642 ? _GEN_158 : _GEN_17; // @[Conditional.scala 39:67]
  assign _GEN_186 = _T_642 ? _GEN_159 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_187 = _T_642 ? _GEN_160 : _GEN_25; // @[Conditional.scala 39:67]
  assign _GEN_188 = _T_642 ? _GEN_161 : _GEN_29; // @[Conditional.scala 39:67]
  assign _GEN_189 = _T_642 ? _GEN_162 : state; // @[Conditional.scala 39:67]
  assign _GEN_190 = _T_588 ? _GEN_109 : active_loop_start_R_control; // @[Conditional.scala 39:67]
  assign _GEN_191 = _T_588 ? _GEN_110 : active_loop_start_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_192 = _T_588 ? _GEN_111 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_193 = _T_588 ? _GEN_112 : active_loop_back_R_control; // @[Conditional.scala 39:67]
  assign _GEN_194 = _T_588 ? _GEN_113 : active_loop_back_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_195 = _T_588 ? _GEN_114 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_196 = _T_588 ? _GEN_115 : _GEN_35; // @[Conditional.scala 39:67]
  assign _GEN_197 = _T_588 ? _GEN_116 : _GEN_37; // @[Conditional.scala 39:67]
  assign _GEN_198 = _T_588 ? _GEN_117 : _GEN_39; // @[Conditional.scala 39:67]
  assign _GEN_199 = _T_588 ? _GEN_118 : _GEN_41; // @[Conditional.scala 39:67]
  assign _GEN_201 = _T_588 ? _GEN_120 : _GEN_34; // @[Conditional.scala 39:67]
  assign _GEN_202 = _T_588 ? _GEN_121 : _GEN_36; // @[Conditional.scala 39:67]
  assign _GEN_203 = _T_588 ? _GEN_122 : _GEN_38; // @[Conditional.scala 39:67]
  assign _GEN_204 = _T_588 ? _GEN_123 : _GEN_40; // @[Conditional.scala 39:67]
  assign _GEN_205 = _T_588 ? _GEN_124 : _GEN_42; // @[Conditional.scala 39:67]
  assign _GEN_206 = _T_588 ? _GEN_125 : _GEN_166; // @[Conditional.scala 39:67]
  assign _GEN_207 = _T_588 ? _GEN_126 : _GEN_167; // @[Conditional.scala 39:67]
  assign _GEN_208 = _T_588 ? _GEN_127 : _GEN_168; // @[Conditional.scala 39:67]
  assign _GEN_209 = _T_588 ? _GEN_128 : _GEN_169; // @[Conditional.scala 39:67]
  assign _GEN_211 = _T_588 ? _GEN_130 : _GEN_171; // @[Conditional.scala 39:67]
  assign _GEN_212 = _T_588 ? _GEN_131 : _GEN_188; // @[Conditional.scala 39:67]
  assign _GEN_213 = _T_588 ? _GEN_132 : _GEN_189; // @[Conditional.scala 39:67]
  assign _GEN_214 = _T_588 ? _GEN_133 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_215 = _T_588 ? _GEN_134 : loop_exit_R_0_control; // @[Conditional.scala 39:67]
  assign _GEN_216 = _T_588 ? _GEN_135 : loop_exit_R_0_taskID; // @[Conditional.scala 39:67]
  assign _GEN_217 = _T_588 ? _GEN_1 : _GEN_163; // @[Conditional.scala 39:67]
  assign _GEN_218 = _T_588 ? _GEN_2 : _GEN_164; // @[Conditional.scala 39:67]
  assign _GEN_219 = _T_588 ? _GEN_3 : _GEN_165; // @[Conditional.scala 39:67]
  assign _GEN_220 = _T_588 ? _GEN_12 : _GEN_172; // @[Conditional.scala 39:67]
  assign _GEN_223 = _T_588 ? _GEN_16 : _GEN_175; // @[Conditional.scala 39:67]
  assign _GEN_224 = _T_588 ? _GEN_15 : _GEN_176; // @[Conditional.scala 39:67]
  assign _GEN_226 = _T_588 ? _GEN_20 : _GEN_178; // @[Conditional.scala 39:67]
  assign _GEN_227 = _T_588 ? _GEN_19 : _GEN_179; // @[Conditional.scala 39:67]
  assign _GEN_229 = _T_588 ? _GEN_24 : _GEN_181; // @[Conditional.scala 39:67]
  assign _GEN_230 = _T_588 ? _GEN_23 : _GEN_182; // @[Conditional.scala 39:67]
  assign _GEN_232 = _T_588 ? _GEN_13 : _GEN_184; // @[Conditional.scala 39:67]
  assign _GEN_233 = _T_588 ? _GEN_17 : _GEN_185; // @[Conditional.scala 39:67]
  assign _GEN_234 = _T_588 ? _GEN_21 : _GEN_186; // @[Conditional.scala 39:67]
  assign _GEN_235 = _T_588 ? _GEN_25 : _GEN_187; // @[Conditional.scala 39:67]
  assign _GEN_236 = _T_565 ? _GEN_59 : _GEN_201; // @[Conditional.scala 40:58]
  assign _GEN_237 = _T_565 ? _GEN_60 : _GEN_202; // @[Conditional.scala 40:58]
  assign _GEN_238 = _T_565 ? _GEN_61 : _GEN_203; // @[Conditional.scala 40:58]
  assign _GEN_239 = _T_565 ? _GEN_62 : _GEN_204; // @[Conditional.scala 40:58]
  assign _GEN_240 = _T_565 ? _GEN_63 : _GEN_205; // @[Conditional.scala 40:58]
  assign _GEN_241 = _T_565 ? _GEN_64 : _GEN_190; // @[Conditional.scala 40:58]
  assign _GEN_242 = _T_565 ? _GEN_65 : _GEN_191; // @[Conditional.scala 40:58]
  assign _GEN_243 = _T_565 ? _GEN_66 : _GEN_192; // @[Conditional.scala 40:58]
  assign _GEN_244 = _T_565 ? _GEN_67 : _GEN_193; // @[Conditional.scala 40:58]
  assign _GEN_245 = _T_565 ? _GEN_68 : _GEN_194; // @[Conditional.scala 40:58]
  assign _GEN_246 = _T_565 ? _GEN_69 : _GEN_195; // @[Conditional.scala 40:58]
  assign _GEN_247 = _T_565 ? _GEN_70 : _GEN_213; // @[Conditional.scala 40:58]
  assign _GEN_248 = _T_565 ? _GEN_71 : _GEN_215; // @[Conditional.scala 40:58]
  assign _GEN_249 = _T_565 ? _GEN_72 : _GEN_216; // @[Conditional.scala 40:58]
  assign _GEN_250 = _T_565 ? _GEN_73 : _GEN_214; // @[Conditional.scala 40:58]
  assign _GEN_251 = _T_565 ? _GEN_35 : _GEN_196; // @[Conditional.scala 40:58]
  assign _GEN_252 = _T_565 ? _GEN_37 : _GEN_197; // @[Conditional.scala 40:58]
  assign _GEN_253 = _T_565 ? _GEN_39 : _GEN_198; // @[Conditional.scala 40:58]
  assign _GEN_254 = _T_565 ? _GEN_41 : _GEN_199; // @[Conditional.scala 40:58]
  assign _GEN_256 = _T_565 ? _GEN_5 : _GEN_206; // @[Conditional.scala 40:58]
  assign _GEN_257 = _T_565 ? _GEN_4 : _GEN_207; // @[Conditional.scala 40:58]
  assign _GEN_258 = _T_565 ? _GEN_6 : _GEN_208; // @[Conditional.scala 40:58]
  assign _GEN_259 = _T_565 ? _GEN_8 : _GEN_209; // @[Conditional.scala 40:58]
  assign _GEN_261 = _T_565 ? _GEN_9 : _GEN_211; // @[Conditional.scala 40:58]
  assign _GEN_262 = _T_565 ? _GEN_29 : _GEN_212; // @[Conditional.scala 40:58]
  assign _GEN_263 = _T_565 ? _GEN_1 : _GEN_217; // @[Conditional.scala 40:58]
  assign _GEN_264 = _T_565 ? _GEN_2 : _GEN_218; // @[Conditional.scala 40:58]
  assign _GEN_265 = _T_565 ? _GEN_3 : _GEN_219; // @[Conditional.scala 40:58]
  assign _GEN_266 = _T_565 ? _GEN_12 : _GEN_220; // @[Conditional.scala 40:58]
  assign _GEN_269 = _T_565 ? _GEN_16 : _GEN_223; // @[Conditional.scala 40:58]
  assign _GEN_270 = _T_565 ? _GEN_15 : _GEN_224; // @[Conditional.scala 40:58]
  assign _GEN_272 = _T_565 ? _GEN_20 : _GEN_226; // @[Conditional.scala 40:58]
  assign _GEN_273 = _T_565 ? _GEN_19 : _GEN_227; // @[Conditional.scala 40:58]
  assign _GEN_275 = _T_565 ? _GEN_24 : _GEN_229; // @[Conditional.scala 40:58]
  assign _GEN_276 = _T_565 ? _GEN_23 : _GEN_230; // @[Conditional.scala 40:58]
  assign _GEN_278 = _T_565 ? _GEN_13 : _GEN_232; // @[Conditional.scala 40:58]
  assign _GEN_279 = _T_565 ? _GEN_17 : _GEN_233; // @[Conditional.scala 40:58]
  assign _GEN_280 = _T_565 ? _GEN_21 : _GEN_234; // @[Conditional.scala 40:58]
  assign _GEN_281 = _T_565 ? _GEN_25 : _GEN_235; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_taskID = in_live_in_R_3_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_taskID = _RAND_13[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_19[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_31[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_34[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_37[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  state = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_519) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_588) begin
          if (_T_519) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_519) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_519) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_519) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_588) begin
          if (_T_519) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_519) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_519) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_519) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_519) begin
            enable_valid_R <= 1'h1;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_519) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_519) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_522) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_522) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_522) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_522) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_522) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_522) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_522) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_522) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_522) begin
          loop_back_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_522) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_522) begin
              loop_back_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_522) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_525) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_525) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_525) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_525) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_8;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_525) begin
          loop_finish_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_525) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_525) begin
              loop_finish_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_525) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_565) begin
        if (_T_528) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_588) begin
          if (_T_528) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_528) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_528) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_531) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_588) begin
          if (_T_531) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_taskID <= 10'h0;
            end else begin
              if (_T_531) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_531) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_565) begin
        if (_T_531) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_588) begin
          if (_T_531) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_531) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_531) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_534) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_588) begin
          if (_T_534) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_taskID <= 10'h0;
            end else begin
              if (_T_534) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_534) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_565) begin
        if (_T_534) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_588) begin
          if (_T_534) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_534) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_534) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_537) begin
          in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
        end
      end else begin
        if (_T_588) begin
          if (_T_537) begin
            in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_taskID <= 10'h0;
            end else begin
              if (_T_537) begin
                in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
              end
            end
          end else begin
            if (_T_537) begin
              in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_565) begin
        if (_T_537) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_588) begin
          if (_T_537) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_537) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_537) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_528) begin
          in_live_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_528) begin
            in_live_in_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_528) begin
                in_live_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_528) begin
              in_live_in_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_531) begin
          in_live_in_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_531) begin
            in_live_in_valid_R_1 <= 1'h1;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              if (_T_531) begin
                in_live_in_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_531) begin
              in_live_in_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_534) begin
          in_live_in_valid_R_2 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_534) begin
            in_live_in_valid_R_2 <= 1'h1;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              if (_T_534) begin
                in_live_in_valid_R_2 <= 1'h1;
              end
            end
          end else begin
            if (_T_534) begin
              in_live_in_valid_R_2 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_537) begin
          in_live_in_valid_R_3 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_537) begin
            in_live_in_valid_R_3 <= 1'h1;
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              if (_T_537) begin
                in_live_in_valid_R_3 <= 1'h1;
              end
            end
          end else begin
            if (_T_537) begin
              in_live_in_valid_R_3 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_540) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_540) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_540) begin
          in_carry_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_540) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_540) begin
              in_carry_in_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_540) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            out_live_in_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_549) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_549) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_549) begin
                out_live_in_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_549) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_0_0 <= _GEN_34;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            out_live_in_valid_R_1_0 <= 1'h1;
          end else begin
            if (_T_552) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_552) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_1_0 <= 1'h1;
            end else begin
              if (_T_552) begin
                out_live_in_valid_R_1_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_552) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_1_0 <= _GEN_36;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            out_live_in_valid_R_2_0 <= 1'h1;
          end else begin
            if (_T_555) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_555) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_2_0 <= 1'h1;
            end else begin
              if (_T_555) begin
                out_live_in_valid_R_2_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_555) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_2_0 <= _GEN_38;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            out_live_in_valid_R_3_0 <= 1'h1;
          end else begin
            if (_T_558) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_558) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_3_0 <= 1'h1;
            end else begin
              if (_T_558) begin
                out_live_in_valid_R_3_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_558) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_3_0 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_549) begin
          out_live_in_fire_R_0_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              if (_T_549) begin
                out_live_in_fire_R_0_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_549) begin
              out_live_in_fire_R_0_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_549) begin
            out_live_in_fire_R_0_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_552) begin
          out_live_in_fire_R_1_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              if (_T_552) begin
                out_live_in_fire_R_1_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_552) begin
              out_live_in_fire_R_1_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_552) begin
            out_live_in_fire_R_1_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_555) begin
          out_live_in_fire_R_2_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              if (_T_555) begin
                out_live_in_fire_R_2_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_555) begin
              out_live_in_fire_R_2_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_555) begin
            out_live_in_fire_R_2_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_558) begin
          out_live_in_fire_R_3_0 <= 1'h1;
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              if (_T_558) begin
                out_live_in_fire_R_3_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_558) begin
              out_live_in_fire_R_3_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_558) begin
            out_live_in_fire_R_3_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            out_carry_out_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_561) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_561) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              out_carry_out_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_561) begin
                out_carry_out_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_561) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_carry_out_valid_R_0_0 <= _GEN_42;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            active_loop_start_R_control <= 1'h1;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            active_loop_start_valid_R <= 1'h1;
          end else begin
            if (_T_542) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_542) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              active_loop_start_valid_R <= 1'h1;
            end else begin
              if (_T_542) begin
                active_loop_start_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_542) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_start_valid_R <= _GEN_30;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_control <= 1'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            active_loop_back_valid_R <= 1'h1;
          end else begin
            if (_T_544) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_544) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              active_loop_back_valid_R <= 1'h1;
            end else begin
              if (_T_544) begin
                active_loop_back_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_544) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_back_valid_R <= _GEN_31;
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 10'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 10'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_control <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_control <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            if (_T_546) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_546) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              if (_T_546) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              if (loop_finish_R_0_control) begin
                loop_exit_valid_R_0 <= 1'h1;
              end else begin
                if (_T_546) begin
                  loop_exit_valid_R_0 <= 1'h0;
                end
              end
            end
          end else begin
            loop_exit_valid_R_0 <= _GEN_32;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_32;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      if (_T_546) begin
        loop_exit_fire_R_0 <= 1'h1;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_565) begin
        if (_T_569) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_588) begin
          if (_T_595) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_642) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [9:0]  io_InLiveIn_0_bits_taskID,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [9:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [9:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [9:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [9:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [9:0]  io_OutLiveIn_field0_0_bits_taskID,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [9:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [9:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [9:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [9:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [9:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [9:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_2;
  reg [9:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_3;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_5;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_6;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_7;
  reg [9:0] in_live_in_R_0_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [9:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [9:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_14;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_15;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_16;
  reg [9:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_17;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_18;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_19;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_20;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_21;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_22;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_23;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_24;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_25;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_26;
  reg [9:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_27;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_28;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_29;
  reg [9:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_30;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_31;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_32;
  reg [9:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_33;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_34;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_35;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_36;
  wire  _T_461; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[LoopBlock.scala 596:26]
  wire  _GEN_2; // @[LoopBlock.scala 596:26]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_464; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_4; // @[LoopBlock.scala 603:33]
  wire  _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_467; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_470; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_12; // @[LoopBlock.scala 623:33]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_473; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_15; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_16; // @[LoopBlock.scala 623:33]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_476; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_19; // @[LoopBlock.scala 623:33]
  wire [31:0] _GEN_20; // @[LoopBlock.scala 623:33]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_479; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_23; // @[LoopBlock.scala 641:37]
  wire [31:0] _GEN_24; // @[LoopBlock.scala 641:37]
  wire  _GEN_25; // @[LoopBlock.scala 641:37]
  wire  _T_481; // @[Decoupled.scala 37:37]
  wire  _GEN_26; // @[LoopBlock.scala 704:39]
  wire  _T_483; // @[Decoupled.scala 37:37]
  wire  _GEN_27; // @[LoopBlock.scala 708:38]
  wire  _T_485; // @[Decoupled.scala 37:37]
  wire  _GEN_28; // @[LoopBlock.scala 713:33]
  wire  _GEN_29; // @[LoopBlock.scala 713:33]
  wire  _T_488; // @[Decoupled.scala 37:37]
  wire  _GEN_30; // @[LoopBlock.scala 722:57]
  wire  _GEN_31; // @[LoopBlock.scala 722:57]
  wire  _T_491; // @[Decoupled.scala 37:37]
  wire  _GEN_32; // @[LoopBlock.scala 722:57]
  wire  _GEN_33; // @[LoopBlock.scala 722:57]
  wire  _T_494; // @[Decoupled.scala 37:37]
  wire  _GEN_34; // @[LoopBlock.scala 722:57]
  wire  _GEN_35; // @[LoopBlock.scala 722:57]
  wire  _T_497; // @[Decoupled.scala 37:37]
  wire  _GEN_36; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_37;
  wire  _T_501; // @[Conditional.scala 37:30]
  wire  _T_502; // @[LoopBlock.scala 765:35]
  wire  _T_503; // @[LoopBlock.scala 765:35]
  wire  _T_504; // @[LoopBlock.scala 869:28]
  wire  _GEN_38; // @[LoopBlock.scala 870:26]
  wire  _GEN_39; // @[LoopBlock.scala 870:26]
  wire  _GEN_40; // @[LoopBlock.scala 870:26]
  wire  _GEN_41; // @[LoopBlock.scala 870:26]
  wire  _GEN_42; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_43; // @[LoopBlock.scala 870:26]
  wire  _GEN_44; // @[LoopBlock.scala 870:26]
  wire  _GEN_45; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_46; // @[LoopBlock.scala 870:26]
  wire  _GEN_47; // @[LoopBlock.scala 870:26]
  wire [1:0] _GEN_48; // @[LoopBlock.scala 870:26]
  wire  _GEN_49; // @[LoopBlock.scala 870:26]
  wire [9:0] _GEN_50; // @[LoopBlock.scala 870:26]
  wire  _GEN_51; // @[LoopBlock.scala 870:26]
  wire  _GEN_52; // @[LoopBlock.scala 869:48]
  wire  _GEN_53; // @[LoopBlock.scala 869:48]
  wire  _GEN_54; // @[LoopBlock.scala 869:48]
  wire  _GEN_55; // @[LoopBlock.scala 869:48]
  wire  _GEN_56; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_57; // @[LoopBlock.scala 869:48]
  wire  _GEN_58; // @[LoopBlock.scala 869:48]
  wire  _GEN_59; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_60; // @[LoopBlock.scala 869:48]
  wire  _GEN_61; // @[LoopBlock.scala 869:48]
  wire [1:0] _GEN_62; // @[LoopBlock.scala 869:48]
  wire  _GEN_63; // @[LoopBlock.scala 869:48]
  wire [9:0] _GEN_64; // @[LoopBlock.scala 869:48]
  wire  _GEN_65; // @[LoopBlock.scala 869:48]
  wire  _T_522; // @[Conditional.scala 37:30]
  wire  _T_523; // @[LoopBlock.scala 898:30]
  wire  _T_526; // @[LoopBlock.scala 828:26]
  wire  _T_527; // @[LoopBlock.scala 828:26]
  wire  _T_528; // @[LoopBlock.scala 899:29]
  wire  _GEN_66; // @[LoopBlock.scala 936:64]
  wire  _GEN_67; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_68; // @[LoopBlock.scala 936:64]
  wire  _GEN_69; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_70; // @[LoopBlock.scala 936:64]
  wire  _GEN_71; // @[LoopBlock.scala 936:64]
  wire [9:0] _GEN_72; // @[LoopBlock.scala 936:64]
  wire [1:0] _GEN_73; // @[LoopBlock.scala 936:64]
  wire  _GEN_74; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_75; // @[LoopBlock.scala 903:56]
  wire  _GEN_76; // @[LoopBlock.scala 903:56]
  wire  _GEN_77; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_78; // @[LoopBlock.scala 903:56]
  wire  _GEN_79; // @[LoopBlock.scala 903:56]
  wire  _GEN_80; // @[LoopBlock.scala 903:56]
  wire  _GEN_81; // @[LoopBlock.scala 903:56]
  wire  _GEN_82; // @[LoopBlock.scala 903:56]
  wire  _GEN_84; // @[LoopBlock.scala 903:56]
  wire  _GEN_85; // @[LoopBlock.scala 903:56]
  wire  _GEN_86; // @[LoopBlock.scala 903:56]
  wire  _GEN_87; // @[LoopBlock.scala 903:56]
  wire  _GEN_88; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_89; // @[LoopBlock.scala 903:56]
  wire  _GEN_90; // @[LoopBlock.scala 903:56]
  wire  _GEN_91; // @[LoopBlock.scala 903:56]
  wire  _GEN_93; // @[LoopBlock.scala 903:56]
  wire  _GEN_94; // @[LoopBlock.scala 903:56]
  wire [1:0] _GEN_95; // @[LoopBlock.scala 903:56]
  wire  _GEN_96; // @[LoopBlock.scala 903:56]
  wire  _GEN_97; // @[LoopBlock.scala 903:56]
  wire [9:0] _GEN_98; // @[LoopBlock.scala 903:56]
  wire  _GEN_99; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_100; // @[LoopBlock.scala 900:55]
  wire  _GEN_101; // @[LoopBlock.scala 900:55]
  wire  _GEN_102; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_103; // @[LoopBlock.scala 900:55]
  wire  _GEN_104; // @[LoopBlock.scala 900:55]
  wire  _GEN_105; // @[LoopBlock.scala 900:55]
  wire  _GEN_106; // @[LoopBlock.scala 900:55]
  wire  _GEN_107; // @[LoopBlock.scala 900:55]
  wire  _GEN_109; // @[LoopBlock.scala 900:55]
  wire  _GEN_110; // @[LoopBlock.scala 900:55]
  wire  _GEN_111; // @[LoopBlock.scala 900:55]
  wire  _GEN_112; // @[LoopBlock.scala 900:55]
  wire  _GEN_113; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_114; // @[LoopBlock.scala 900:55]
  wire  _GEN_115; // @[LoopBlock.scala 900:55]
  wire  _GEN_116; // @[LoopBlock.scala 900:55]
  wire  _GEN_118; // @[LoopBlock.scala 900:55]
  wire  _GEN_119; // @[LoopBlock.scala 900:55]
  wire [1:0] _GEN_120; // @[LoopBlock.scala 900:55]
  wire  _GEN_121; // @[LoopBlock.scala 900:55]
  wire  _GEN_122; // @[LoopBlock.scala 900:55]
  wire [9:0] _GEN_123; // @[LoopBlock.scala 900:55]
  wire  _T_573; // @[Conditional.scala 37:30]
  wire [9:0] _GEN_124; // @[LoopBlock.scala 955:48]
  wire  _GEN_125; // @[LoopBlock.scala 955:48]
  wire  _GEN_126; // @[LoopBlock.scala 955:48]
  wire  _GEN_127; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_128; // @[LoopBlock.scala 955:48]
  wire  _GEN_129; // @[LoopBlock.scala 955:48]
  wire  _GEN_130; // @[LoopBlock.scala 955:48]
  wire  _GEN_132; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_133; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_134; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_136; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_137; // @[LoopBlock.scala 955:48]
  wire [31:0] _GEN_139; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_140; // @[LoopBlock.scala 955:48]
  wire  _GEN_142; // @[LoopBlock.scala 955:48]
  wire  _GEN_143; // @[LoopBlock.scala 955:48]
  wire  _GEN_144; // @[LoopBlock.scala 955:48]
  wire  _GEN_145; // @[LoopBlock.scala 955:48]
  wire [1:0] _GEN_146; // @[LoopBlock.scala 955:48]
  wire [9:0] _GEN_147; // @[Conditional.scala 39:67]
  wire  _GEN_148; // @[Conditional.scala 39:67]
  wire  _GEN_149; // @[Conditional.scala 39:67]
  wire  _GEN_150; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_151; // @[Conditional.scala 39:67]
  wire  _GEN_152; // @[Conditional.scala 39:67]
  wire  _GEN_153; // @[Conditional.scala 39:67]
  wire  _GEN_155; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_156; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_157; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_159; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_160; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_162; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_163; // @[Conditional.scala 39:67]
  wire  _GEN_165; // @[Conditional.scala 39:67]
  wire  _GEN_166; // @[Conditional.scala 39:67]
  wire  _GEN_167; // @[Conditional.scala 39:67]
  wire  _GEN_168; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_169; // @[Conditional.scala 39:67]
  wire  _GEN_170; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_171; // @[Conditional.scala 39:67]
  wire  _GEN_172; // @[Conditional.scala 39:67]
  wire  _GEN_173; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_174; // @[Conditional.scala 39:67]
  wire  _GEN_175; // @[Conditional.scala 39:67]
  wire  _GEN_176; // @[Conditional.scala 39:67]
  wire  _GEN_177; // @[Conditional.scala 39:67]
  wire  _GEN_178; // @[Conditional.scala 39:67]
  wire  _GEN_180; // @[Conditional.scala 39:67]
  wire  _GEN_181; // @[Conditional.scala 39:67]
  wire  _GEN_182; // @[Conditional.scala 39:67]
  wire  _GEN_183; // @[Conditional.scala 39:67]
  wire  _GEN_184; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_185; // @[Conditional.scala 39:67]
  wire  _GEN_186; // @[Conditional.scala 39:67]
  wire  _GEN_187; // @[Conditional.scala 39:67]
  wire  _GEN_189; // @[Conditional.scala 39:67]
  wire  _GEN_190; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_191; // @[Conditional.scala 39:67]
  wire  _GEN_192; // @[Conditional.scala 39:67]
  wire  _GEN_193; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_194; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_195; // @[Conditional.scala 39:67]
  wire  _GEN_196; // @[Conditional.scala 39:67]
  wire  _GEN_197; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_198; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_199; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_201; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_202; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_204; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_205; // @[Conditional.scala 39:67]
  wire  _GEN_207; // @[Conditional.scala 39:67]
  wire  _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_209; // @[Conditional.scala 39:67]
  wire  _GEN_210; // @[Conditional.scala 40:58]
  wire  _GEN_211; // @[Conditional.scala 40:58]
  wire  _GEN_212; // @[Conditional.scala 40:58]
  wire  _GEN_213; // @[Conditional.scala 40:58]
  wire  _GEN_214; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_215; // @[Conditional.scala 40:58]
  wire  _GEN_216; // @[Conditional.scala 40:58]
  wire  _GEN_217; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_218; // @[Conditional.scala 40:58]
  wire  _GEN_219; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_220; // @[Conditional.scala 40:58]
  wire  _GEN_221; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_222; // @[Conditional.scala 40:58]
  wire  _GEN_223; // @[Conditional.scala 40:58]
  wire  _GEN_224; // @[Conditional.scala 40:58]
  wire  _GEN_225; // @[Conditional.scala 40:58]
  wire  _GEN_226; // @[Conditional.scala 40:58]
  wire  _GEN_228; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_229; // @[Conditional.scala 40:58]
  wire  _GEN_230; // @[Conditional.scala 40:58]
  wire  _GEN_231; // @[Conditional.scala 40:58]
  wire  _GEN_233; // @[Conditional.scala 40:58]
  wire  _GEN_234; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_235; // @[Conditional.scala 40:58]
  wire  _GEN_236; // @[Conditional.scala 40:58]
  wire  _GEN_237; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_238; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_239; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_241; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_242; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_244; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_245; // @[Conditional.scala 40:58]
  wire  _GEN_247; // @[Conditional.scala 40:58]
  wire  _GEN_248; // @[Conditional.scala 40:58]
  wire  _GEN_249; // @[Conditional.scala 40:58]
  assign _T_461 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_461 ? io_enable_bits_taskID : enable_R_taskID; // @[LoopBlock.scala 596:26]
  assign _GEN_2 = _T_461 ? io_enable_bits_control : enable_R_control; // @[LoopBlock.scala 596:26]
  assign _GEN_3 = _T_461 ? 1'h1 : enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_464 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_464 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_464 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_464 ? 1'h1 : loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_467 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_467 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_467 ? 1'h1 : loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_470 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_470 ? io_InLiveIn_0_bits_taskID : in_live_in_R_0_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_12 = _T_470 ? io_InLiveIn_0_bits_data : in_live_in_R_0_data; // @[LoopBlock.scala 623:33]
  assign _GEN_13 = _T_470 ? 1'h1 : in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_473 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_15 = _T_473 ? io_InLiveIn_1_bits_taskID : in_live_in_R_1_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_16 = _T_473 ? io_InLiveIn_1_bits_data : in_live_in_R_1_data; // @[LoopBlock.scala 623:33]
  assign _GEN_17 = _T_473 ? 1'h1 : in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_476 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_19 = _T_476 ? io_InLiveIn_2_bits_taskID : in_live_in_R_2_taskID; // @[LoopBlock.scala 623:33]
  assign _GEN_20 = _T_476 ? io_InLiveIn_2_bits_data : in_live_in_R_2_data; // @[LoopBlock.scala 623:33]
  assign _GEN_21 = _T_476 ? 1'h1 : in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_479 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_23 = _T_479 ? io_CarryDepenIn_0_bits_taskID : in_carry_in_R_0_taskID; // @[LoopBlock.scala 641:37]
  assign _GEN_24 = _T_479 ? io_CarryDepenIn_0_bits_data : in_carry_in_R_0_data; // @[LoopBlock.scala 641:37]
  assign _GEN_25 = _T_479 ? 1'h1 : in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_481 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 37:37]
  assign _GEN_26 = _T_481 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_483 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 37:37]
  assign _GEN_27 = _T_483 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_485 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_28 = _T_485 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_29 = _T_485 ? 1'h1 : loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_488 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_30 = _T_488 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_31 = _T_488 ? 1'h1 : out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_491 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_32 = _T_491 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_33 = _T_491 ? 1'h1 : out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_494 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_34 = _T_494 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_35 = _T_494 ? 1'h1 : out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_497 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_36 = _T_497 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_501 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_502 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_503 = _T_502 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_504 = _T_503 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_38 = enable_R_control ? 1'h1 : _GEN_30; // @[LoopBlock.scala 870:26]
  assign _GEN_39 = enable_R_control ? 1'h1 : _GEN_32; // @[LoopBlock.scala 870:26]
  assign _GEN_40 = enable_R_control ? 1'h1 : _GEN_34; // @[LoopBlock.scala 870:26]
  assign _GEN_41 = enable_R_control ? 1'h1 : _GEN_36; // @[LoopBlock.scala 870:26]
  assign _GEN_42 = enable_R_control ? 1'h1 : active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_43 = enable_R_control ? enable_R_taskID : active_loop_start_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_44 = enable_R_control ? 1'h1 : _GEN_26; // @[LoopBlock.scala 870:26]
  assign _GEN_45 = enable_R_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_46 = enable_R_control ? enable_R_taskID : active_loop_back_R_taskID; // @[LoopBlock.scala 870:26]
  assign _GEN_47 = enable_R_control ? 1'h1 : _GEN_27; // @[LoopBlock.scala 870:26]
  assign _GEN_48 = enable_R_control ? 2'h1 : 2'h2; // @[LoopBlock.scala 870:26]
  assign _GEN_49 = enable_R_control ? loop_exit_R_0_control : 1'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_50 = enable_R_control ? loop_exit_R_0_taskID : 10'h0; // @[LoopBlock.scala 870:26]
  assign _GEN_51 = enable_R_control ? _GEN_28 : 1'h1; // @[LoopBlock.scala 870:26]
  assign _GEN_52 = _T_504 ? _GEN_38 : _GEN_30; // @[LoopBlock.scala 869:48]
  assign _GEN_53 = _T_504 ? _GEN_39 : _GEN_32; // @[LoopBlock.scala 869:48]
  assign _GEN_54 = _T_504 ? _GEN_40 : _GEN_34; // @[LoopBlock.scala 869:48]
  assign _GEN_55 = _T_504 ? _GEN_41 : _GEN_36; // @[LoopBlock.scala 869:48]
  assign _GEN_56 = _T_504 ? _GEN_42 : active_loop_start_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_57 = _T_504 ? _GEN_43 : active_loop_start_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_58 = _T_504 ? _GEN_44 : _GEN_26; // @[LoopBlock.scala 869:48]
  assign _GEN_59 = _T_504 ? _GEN_45 : active_loop_back_R_control; // @[LoopBlock.scala 869:48]
  assign _GEN_60 = _T_504 ? _GEN_46 : active_loop_back_R_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_61 = _T_504 ? _GEN_47 : _GEN_27; // @[LoopBlock.scala 869:48]
  assign _GEN_62 = _T_504 ? _GEN_48 : state; // @[LoopBlock.scala 869:48]
  assign _GEN_63 = _T_504 ? _GEN_49 : loop_exit_R_0_control; // @[LoopBlock.scala 869:48]
  assign _GEN_64 = _T_504 ? _GEN_50 : loop_exit_R_0_taskID; // @[LoopBlock.scala 869:48]
  assign _GEN_65 = _T_504 ? _GEN_51 : _GEN_28; // @[LoopBlock.scala 869:48]
  assign _T_522 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_523 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_526 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_527 = _T_526 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_528 = _T_523 & _T_527; // @[LoopBlock.scala 899:29]
  assign _GEN_66 = loop_finish_R_0_control ? 1'h1 : _GEN_28; // @[LoopBlock.scala 936:64]
  assign _GEN_67 = loop_finish_R_0_control ? 1'h0 : active_loop_start_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_68 = loop_finish_R_0_control ? 10'h0 : active_loop_start_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_69 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_70 = loop_finish_R_0_control ? 10'h0 : active_loop_back_R_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_71 = loop_finish_R_0_control ? 1'h1 : loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_72 = loop_finish_R_0_control ? loop_back_R_0_taskID : loop_exit_R_0_taskID; // @[LoopBlock.scala 936:64]
  assign _GEN_73 = loop_finish_R_0_control ? 2'h2 : state; // @[LoopBlock.scala 936:64]
  assign _GEN_74 = loop_back_R_0_control ? 1'h0 : _GEN_67; // @[LoopBlock.scala 903:56]
  assign _GEN_75 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_68; // @[LoopBlock.scala 903:56]
  assign _GEN_76 = loop_back_R_0_control ? 1'h1 : _GEN_26; // @[LoopBlock.scala 903:56]
  assign _GEN_77 = loop_back_R_0_control ? 1'h1 : _GEN_69; // @[LoopBlock.scala 903:56]
  assign _GEN_78 = loop_back_R_0_control ? loop_back_R_0_taskID : _GEN_70; // @[LoopBlock.scala 903:56]
  assign _GEN_79 = loop_back_R_0_control ? 1'h1 : _GEN_27; // @[LoopBlock.scala 903:56]
  assign _GEN_80 = loop_back_R_0_control ? 1'h0 : _GEN_31; // @[LoopBlock.scala 903:56]
  assign _GEN_81 = loop_back_R_0_control ? 1'h0 : _GEN_33; // @[LoopBlock.scala 903:56]
  assign _GEN_82 = loop_back_R_0_control ? 1'h0 : _GEN_35; // @[LoopBlock.scala 903:56]
  assign _GEN_84 = loop_back_R_0_control ? 1'h1 : _GEN_30; // @[LoopBlock.scala 903:56]
  assign _GEN_85 = loop_back_R_0_control ? 1'h1 : _GEN_32; // @[LoopBlock.scala 903:56]
  assign _GEN_86 = loop_back_R_0_control ? 1'h1 : _GEN_34; // @[LoopBlock.scala 903:56]
  assign _GEN_87 = loop_back_R_0_control ? 1'h1 : _GEN_36; // @[LoopBlock.scala 903:56]
  assign _GEN_88 = loop_back_R_0_control ? 1'h0 : _GEN_5; // @[LoopBlock.scala 903:56]
  assign _GEN_89 = loop_back_R_0_control ? 10'h0 : _GEN_4; // @[LoopBlock.scala 903:56]
  assign _GEN_90 = loop_back_R_0_control ? 1'h0 : _GEN_6; // @[LoopBlock.scala 903:56]
  assign _GEN_91 = loop_back_R_0_control ? 1'h0 : _GEN_8; // @[LoopBlock.scala 903:56]
  assign _GEN_93 = loop_back_R_0_control ? 1'h0 : _GEN_9; // @[LoopBlock.scala 903:56]
  assign _GEN_94 = loop_back_R_0_control ? 1'h0 : _GEN_25; // @[LoopBlock.scala 903:56]
  assign _GEN_95 = loop_back_R_0_control ? 2'h1 : _GEN_73; // @[LoopBlock.scala 903:56]
  assign _GEN_96 = loop_back_R_0_control ? _GEN_28 : _GEN_66; // @[LoopBlock.scala 903:56]
  assign _GEN_97 = loop_back_R_0_control ? loop_exit_R_0_control : _GEN_71; // @[LoopBlock.scala 903:56]
  assign _GEN_98 = loop_back_R_0_control ? loop_exit_R_0_taskID : _GEN_72; // @[LoopBlock.scala 903:56]
  assign _GEN_99 = _T_528 ? _GEN_74 : active_loop_start_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_100 = _T_528 ? _GEN_75 : active_loop_start_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_101 = _T_528 ? _GEN_76 : _GEN_26; // @[LoopBlock.scala 900:55]
  assign _GEN_102 = _T_528 ? _GEN_77 : active_loop_back_R_control; // @[LoopBlock.scala 900:55]
  assign _GEN_103 = _T_528 ? _GEN_78 : active_loop_back_R_taskID; // @[LoopBlock.scala 900:55]
  assign _GEN_104 = _T_528 ? _GEN_79 : _GEN_27; // @[LoopBlock.scala 900:55]
  assign _GEN_105 = _T_528 ? _GEN_80 : _GEN_31; // @[LoopBlock.scala 900:55]
  assign _GEN_106 = _T_528 ? _GEN_81 : _GEN_33; // @[LoopBlock.scala 900:55]
  assign _GEN_107 = _T_528 ? _GEN_82 : _GEN_35; // @[LoopBlock.scala 900:55]
  assign _GEN_109 = _T_528 ? _GEN_84 : _GEN_30; // @[LoopBlock.scala 900:55]
  assign _GEN_110 = _T_528 ? _GEN_85 : _GEN_32; // @[LoopBlock.scala 900:55]
  assign _GEN_111 = _T_528 ? _GEN_86 : _GEN_34; // @[LoopBlock.scala 900:55]
  assign _GEN_112 = _T_528 ? _GEN_87 : _GEN_36; // @[LoopBlock.scala 900:55]
  assign _GEN_113 = _T_528 ? _GEN_88 : _GEN_5; // @[LoopBlock.scala 900:55]
  assign _GEN_114 = _T_528 ? _GEN_89 : _GEN_4; // @[LoopBlock.scala 900:55]
  assign _GEN_115 = _T_528 ? _GEN_90 : _GEN_6; // @[LoopBlock.scala 900:55]
  assign _GEN_116 = _T_528 ? _GEN_91 : _GEN_8; // @[LoopBlock.scala 900:55]
  assign _GEN_118 = _T_528 ? _GEN_93 : _GEN_9; // @[LoopBlock.scala 900:55]
  assign _GEN_119 = _T_528 ? _GEN_94 : _GEN_25; // @[LoopBlock.scala 900:55]
  assign _GEN_120 = _T_528 ? _GEN_95 : state; // @[LoopBlock.scala 900:55]
  assign _GEN_121 = _T_528 ? _GEN_96 : _GEN_28; // @[LoopBlock.scala 900:55]
  assign _GEN_122 = _T_528 ? _GEN_97 : loop_exit_R_0_control; // @[LoopBlock.scala 900:55]
  assign _GEN_123 = _T_528 ? _GEN_98 : loop_exit_R_0_taskID; // @[LoopBlock.scala 900:55]
  assign _T_573 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_124 = loop_exit_fire_R_0 ? 10'h0 : _GEN_1; // @[LoopBlock.scala 955:48]
  assign _GEN_125 = loop_exit_fire_R_0 ? 1'h0 : _GEN_2; // @[LoopBlock.scala 955:48]
  assign _GEN_126 = loop_exit_fire_R_0 ? 1'h0 : _GEN_3; // @[LoopBlock.scala 955:48]
  assign _GEN_127 = loop_exit_fire_R_0 ? 1'h0 : _GEN_5; // @[LoopBlock.scala 955:48]
  assign _GEN_128 = loop_exit_fire_R_0 ? 10'h0 : _GEN_4; // @[LoopBlock.scala 955:48]
  assign _GEN_129 = loop_exit_fire_R_0 ? 1'h0 : _GEN_6; // @[LoopBlock.scala 955:48]
  assign _GEN_130 = loop_exit_fire_R_0 ? 1'h0 : _GEN_8; // @[LoopBlock.scala 955:48]
  assign _GEN_132 = loop_exit_fire_R_0 ? 1'h0 : _GEN_9; // @[LoopBlock.scala 955:48]
  assign _GEN_133 = loop_exit_fire_R_0 ? 32'h0 : _GEN_12; // @[LoopBlock.scala 955:48]
  assign _GEN_134 = loop_exit_fire_R_0 ? 10'h0 : _GEN_11; // @[LoopBlock.scala 955:48]
  assign _GEN_136 = loop_exit_fire_R_0 ? 32'h0 : _GEN_16; // @[LoopBlock.scala 955:48]
  assign _GEN_137 = loop_exit_fire_R_0 ? 10'h0 : _GEN_15; // @[LoopBlock.scala 955:48]
  assign _GEN_139 = loop_exit_fire_R_0 ? 32'h0 : _GEN_20; // @[LoopBlock.scala 955:48]
  assign _GEN_140 = loop_exit_fire_R_0 ? 10'h0 : _GEN_19; // @[LoopBlock.scala 955:48]
  assign _GEN_142 = loop_exit_fire_R_0 ? 1'h0 : _GEN_13; // @[LoopBlock.scala 955:48]
  assign _GEN_143 = loop_exit_fire_R_0 ? 1'h0 : _GEN_17; // @[LoopBlock.scala 955:48]
  assign _GEN_144 = loop_exit_fire_R_0 ? 1'h0 : _GEN_21; // @[LoopBlock.scala 955:48]
  assign _GEN_145 = loop_exit_fire_R_0 ? 1'h0 : _GEN_25; // @[LoopBlock.scala 955:48]
  assign _GEN_146 = loop_exit_fire_R_0 ? 2'h0 : state; // @[LoopBlock.scala 955:48]
  assign _GEN_147 = _T_573 ? _GEN_124 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_148 = _T_573 ? _GEN_125 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_149 = _T_573 ? _GEN_126 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_150 = _T_573 ? _GEN_127 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_151 = _T_573 ? _GEN_128 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_152 = _T_573 ? _GEN_129 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_153 = _T_573 ? _GEN_130 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_155 = _T_573 ? _GEN_132 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_156 = _T_573 ? _GEN_133 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_157 = _T_573 ? _GEN_134 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_159 = _T_573 ? _GEN_136 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_160 = _T_573 ? _GEN_137 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_162 = _T_573 ? _GEN_139 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_163 = _T_573 ? _GEN_140 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_165 = _T_573 ? _GEN_142 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_166 = _T_573 ? _GEN_143 : _GEN_17; // @[Conditional.scala 39:67]
  assign _GEN_167 = _T_573 ? _GEN_144 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_168 = _T_573 ? _GEN_145 : _GEN_25; // @[Conditional.scala 39:67]
  assign _GEN_169 = _T_573 ? _GEN_146 : state; // @[Conditional.scala 39:67]
  assign _GEN_170 = _T_522 ? _GEN_99 : active_loop_start_R_control; // @[Conditional.scala 39:67]
  assign _GEN_171 = _T_522 ? _GEN_100 : active_loop_start_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_172 = _T_522 ? _GEN_101 : _GEN_26; // @[Conditional.scala 39:67]
  assign _GEN_173 = _T_522 ? _GEN_102 : active_loop_back_R_control; // @[Conditional.scala 39:67]
  assign _GEN_174 = _T_522 ? _GEN_103 : active_loop_back_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_175 = _T_522 ? _GEN_104 : _GEN_27; // @[Conditional.scala 39:67]
  assign _GEN_176 = _T_522 ? _GEN_105 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_177 = _T_522 ? _GEN_106 : _GEN_33; // @[Conditional.scala 39:67]
  assign _GEN_178 = _T_522 ? _GEN_107 : _GEN_35; // @[Conditional.scala 39:67]
  assign _GEN_180 = _T_522 ? _GEN_109 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_181 = _T_522 ? _GEN_110 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_182 = _T_522 ? _GEN_111 : _GEN_34; // @[Conditional.scala 39:67]
  assign _GEN_183 = _T_522 ? _GEN_112 : _GEN_36; // @[Conditional.scala 39:67]
  assign _GEN_184 = _T_522 ? _GEN_113 : _GEN_150; // @[Conditional.scala 39:67]
  assign _GEN_185 = _T_522 ? _GEN_114 : _GEN_151; // @[Conditional.scala 39:67]
  assign _GEN_186 = _T_522 ? _GEN_115 : _GEN_152; // @[Conditional.scala 39:67]
  assign _GEN_187 = _T_522 ? _GEN_116 : _GEN_153; // @[Conditional.scala 39:67]
  assign _GEN_189 = _T_522 ? _GEN_118 : _GEN_155; // @[Conditional.scala 39:67]
  assign _GEN_190 = _T_522 ? _GEN_119 : _GEN_168; // @[Conditional.scala 39:67]
  assign _GEN_191 = _T_522 ? _GEN_120 : _GEN_169; // @[Conditional.scala 39:67]
  assign _GEN_192 = _T_522 ? _GEN_121 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_193 = _T_522 ? _GEN_122 : loop_exit_R_0_control; // @[Conditional.scala 39:67]
  assign _GEN_194 = _T_522 ? _GEN_123 : loop_exit_R_0_taskID; // @[Conditional.scala 39:67]
  assign _GEN_195 = _T_522 ? _GEN_1 : _GEN_147; // @[Conditional.scala 39:67]
  assign _GEN_196 = _T_522 ? _GEN_2 : _GEN_148; // @[Conditional.scala 39:67]
  assign _GEN_197 = _T_522 ? _GEN_3 : _GEN_149; // @[Conditional.scala 39:67]
  assign _GEN_198 = _T_522 ? _GEN_12 : _GEN_156; // @[Conditional.scala 39:67]
  assign _GEN_199 = _T_522 ? _GEN_11 : _GEN_157; // @[Conditional.scala 39:67]
  assign _GEN_201 = _T_522 ? _GEN_16 : _GEN_159; // @[Conditional.scala 39:67]
  assign _GEN_202 = _T_522 ? _GEN_15 : _GEN_160; // @[Conditional.scala 39:67]
  assign _GEN_204 = _T_522 ? _GEN_20 : _GEN_162; // @[Conditional.scala 39:67]
  assign _GEN_205 = _T_522 ? _GEN_19 : _GEN_163; // @[Conditional.scala 39:67]
  assign _GEN_207 = _T_522 ? _GEN_13 : _GEN_165; // @[Conditional.scala 39:67]
  assign _GEN_208 = _T_522 ? _GEN_17 : _GEN_166; // @[Conditional.scala 39:67]
  assign _GEN_209 = _T_522 ? _GEN_21 : _GEN_167; // @[Conditional.scala 39:67]
  assign _GEN_210 = _T_501 ? _GEN_52 : _GEN_180; // @[Conditional.scala 40:58]
  assign _GEN_211 = _T_501 ? _GEN_53 : _GEN_181; // @[Conditional.scala 40:58]
  assign _GEN_212 = _T_501 ? _GEN_54 : _GEN_182; // @[Conditional.scala 40:58]
  assign _GEN_213 = _T_501 ? _GEN_55 : _GEN_183; // @[Conditional.scala 40:58]
  assign _GEN_214 = _T_501 ? _GEN_56 : _GEN_170; // @[Conditional.scala 40:58]
  assign _GEN_215 = _T_501 ? _GEN_57 : _GEN_171; // @[Conditional.scala 40:58]
  assign _GEN_216 = _T_501 ? _GEN_58 : _GEN_172; // @[Conditional.scala 40:58]
  assign _GEN_217 = _T_501 ? _GEN_59 : _GEN_173; // @[Conditional.scala 40:58]
  assign _GEN_218 = _T_501 ? _GEN_60 : _GEN_174; // @[Conditional.scala 40:58]
  assign _GEN_219 = _T_501 ? _GEN_61 : _GEN_175; // @[Conditional.scala 40:58]
  assign _GEN_220 = _T_501 ? _GEN_62 : _GEN_191; // @[Conditional.scala 40:58]
  assign _GEN_221 = _T_501 ? _GEN_63 : _GEN_193; // @[Conditional.scala 40:58]
  assign _GEN_222 = _T_501 ? _GEN_64 : _GEN_194; // @[Conditional.scala 40:58]
  assign _GEN_223 = _T_501 ? _GEN_65 : _GEN_192; // @[Conditional.scala 40:58]
  assign _GEN_224 = _T_501 ? _GEN_31 : _GEN_176; // @[Conditional.scala 40:58]
  assign _GEN_225 = _T_501 ? _GEN_33 : _GEN_177; // @[Conditional.scala 40:58]
  assign _GEN_226 = _T_501 ? _GEN_35 : _GEN_178; // @[Conditional.scala 40:58]
  assign _GEN_228 = _T_501 ? _GEN_5 : _GEN_184; // @[Conditional.scala 40:58]
  assign _GEN_229 = _T_501 ? _GEN_4 : _GEN_185; // @[Conditional.scala 40:58]
  assign _GEN_230 = _T_501 ? _GEN_6 : _GEN_186; // @[Conditional.scala 40:58]
  assign _GEN_231 = _T_501 ? _GEN_8 : _GEN_187; // @[Conditional.scala 40:58]
  assign _GEN_233 = _T_501 ? _GEN_9 : _GEN_189; // @[Conditional.scala 40:58]
  assign _GEN_234 = _T_501 ? _GEN_25 : _GEN_190; // @[Conditional.scala 40:58]
  assign _GEN_235 = _T_501 ? _GEN_1 : _GEN_195; // @[Conditional.scala 40:58]
  assign _GEN_236 = _T_501 ? _GEN_2 : _GEN_196; // @[Conditional.scala 40:58]
  assign _GEN_237 = _T_501 ? _GEN_3 : _GEN_197; // @[Conditional.scala 40:58]
  assign _GEN_238 = _T_501 ? _GEN_12 : _GEN_198; // @[Conditional.scala 40:58]
  assign _GEN_239 = _T_501 ? _GEN_11 : _GEN_199; // @[Conditional.scala 40:58]
  assign _GEN_241 = _T_501 ? _GEN_16 : _GEN_201; // @[Conditional.scala 40:58]
  assign _GEN_242 = _T_501 ? _GEN_15 : _GEN_202; // @[Conditional.scala 40:58]
  assign _GEN_244 = _T_501 ? _GEN_20 : _GEN_204; // @[Conditional.scala 40:58]
  assign _GEN_245 = _T_501 ? _GEN_19 : _GEN_205; // @[Conditional.scala 40:58]
  assign _GEN_247 = _T_501 ? _GEN_13 : _GEN_207; // @[Conditional.scala 40:58]
  assign _GEN_248 = _T_501 ? _GEN_17 : _GEN_208; // @[Conditional.scala 40:58]
  assign _GEN_249 = _T_501 ? _GEN_21 : _GEN_209; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_taskID = in_live_in_R_0_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  in_live_in_R_0_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_27[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_30[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_33[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  state = _RAND_37[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_461) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_522) begin
          if (_T_461) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_461) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_461) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_461) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_522) begin
          if (_T_461) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_461) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_461) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_461) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_461) begin
            enable_valid_R <= 1'h1;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_461) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_461) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_464) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_464) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_464) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 10'h0;
            end else begin
              if (_T_464) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_464) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_464) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_464) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_464) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_464) begin
          loop_back_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_464) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_464) begin
              loop_back_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              if (_T_464) begin
                loop_back_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_467) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_467) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_467) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_467) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_8;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_467) begin
          loop_finish_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_467) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_467) begin
              loop_finish_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              if (_T_467) begin
                loop_finish_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_470) begin
          in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
        end
      end else begin
        if (_T_522) begin
          if (_T_470) begin
            in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_taskID <= 10'h0;
            end else begin
              if (_T_470) begin
                in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
              end
            end
          end else begin
            if (_T_470) begin
              in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_501) begin
        if (_T_470) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_522) begin
          if (_T_470) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_470) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_470) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_473) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_522) begin
          if (_T_473) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_taskID <= 10'h0;
            end else begin
              if (_T_473) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_473) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_501) begin
        if (_T_473) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_522) begin
          if (_T_473) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_473) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_473) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_476) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_522) begin
          if (_T_476) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_taskID <= 10'h0;
            end else begin
              if (_T_476) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_476) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_501) begin
        if (_T_476) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_522) begin
          if (_T_476) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_476) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_476) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_470) begin
          in_live_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_470) begin
            in_live_in_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_470) begin
                in_live_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_470) begin
              in_live_in_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_473) begin
          in_live_in_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_473) begin
            in_live_in_valid_R_1 <= 1'h1;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              if (_T_473) begin
                in_live_in_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_473) begin
              in_live_in_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_476) begin
          in_live_in_valid_R_2 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_476) begin
            in_live_in_valid_R_2 <= 1'h1;
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              if (_T_476) begin
                in_live_in_valid_R_2 <= 1'h1;
              end
            end
          end else begin
            if (_T_476) begin
              in_live_in_valid_R_2 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_479) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_479) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_479) begin
          in_carry_in_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_479) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_479) begin
              in_carry_in_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              if (_T_479) begin
                in_carry_in_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            out_live_in_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_488) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_488) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_488) begin
                out_live_in_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_488) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_0_0 <= _GEN_30;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            out_live_in_valid_R_1_0 <= 1'h1;
          end else begin
            if (_T_491) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_491) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_1_0 <= 1'h1;
            end else begin
              if (_T_491) begin
                out_live_in_valid_R_1_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_491) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_1_0 <= _GEN_32;
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            out_live_in_valid_R_2_0 <= 1'h1;
          end else begin
            if (_T_494) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_494) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_live_in_valid_R_2_0 <= 1'h1;
            end else begin
              if (_T_494) begin
                out_live_in_valid_R_2_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_494) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          out_live_in_valid_R_2_0 <= _GEN_34;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_488) begin
          out_live_in_fire_R_0_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              if (_T_488) begin
                out_live_in_fire_R_0_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_488) begin
              out_live_in_fire_R_0_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_488) begin
            out_live_in_fire_R_0_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_491) begin
          out_live_in_fire_R_1_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              if (_T_491) begin
                out_live_in_fire_R_1_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_491) begin
              out_live_in_fire_R_1_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_491) begin
            out_live_in_fire_R_1_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_494) begin
          out_live_in_fire_R_2_0 <= 1'h1;
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              if (_T_494) begin
                out_live_in_fire_R_2_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_494) begin
              out_live_in_fire_R_2_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_494) begin
            out_live_in_fire_R_2_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            out_carry_out_valid_R_0_0 <= 1'h1;
          end else begin
            if (_T_497) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_497) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              out_carry_out_valid_R_0_0 <= 1'h1;
            end else begin
              if (_T_497) begin
                out_carry_out_valid_R_0_0 <= 1'h0;
              end
            end
          end else begin
            if (_T_497) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_carry_out_valid_R_0_0 <= _GEN_36;
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            active_loop_start_R_control <= 1'h1;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            active_loop_start_valid_R <= 1'h1;
          end else begin
            if (_T_481) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_481) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              active_loop_start_valid_R <= 1'h1;
            end else begin
              if (_T_481) begin
                active_loop_start_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_481) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_start_valid_R <= _GEN_26;
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 10'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_control <= 1'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            active_loop_back_valid_R <= 1'h1;
          end else begin
            if (_T_483) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_483) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              active_loop_back_valid_R <= 1'h1;
            end else begin
              if (_T_483) begin
                active_loop_back_valid_R <= 1'h0;
              end
            end
          end else begin
            if (_T_483) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          active_loop_back_valid_R <= _GEN_27;
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 10'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 10'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_control <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_control <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            if (_T_485) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_485) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              if (_T_485) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              if (loop_finish_R_0_control) begin
                loop_exit_valid_R_0 <= 1'h1;
              end else begin
                if (_T_485) begin
                  loop_exit_valid_R_0 <= 1'h0;
                end
              end
            end
          end else begin
            loop_exit_valid_R_0 <= _GEN_28;
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_28;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      if (_T_485) begin
        loop_exit_fire_R_0 <= 1'h1;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_501) begin
        if (_T_504) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_522) begin
          if (_T_528) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_573) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module BasicBlockNoMaskFastNode(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [9:0] in_data_R_0_taskID; // @[BasicBlock.scala 988:46]
  reg [31:0] _RAND_0;
  reg  in_data_R_0_control; // @[BasicBlock.scala 988:46]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 989:52]
  reg [31:0] _RAND_2;
  reg [9:0] output_R_taskID; // @[BasicBlock.scala 991:25]
  reg [31:0] _RAND_3;
  reg  output_R_control; // @[BasicBlock.scala 991:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 992:49]
  reg [31:0] _RAND_5;
  reg  output_fire_R_0; // @[BasicBlock.scala 993:48]
  reg [31:0] _RAND_6;
  wire  _T_73; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[BasicBlock.scala 998:36]
  wire  _GEN_2; // @[BasicBlock.scala 998:36]
  wire  _GEN_3; // @[BasicBlock.scala 998:36]
  wire [9:0] in_task_ID; // @[BasicBlock.scala 1005:34]
  wire  _T_75; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[BasicBlock.scala 1010:28]
  wire  _GEN_5; // @[BasicBlock.scala 1010:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 1027:85]
  reg  state; // @[BasicBlock.scala 1040:22]
  reg [31:0] _RAND_7;
  wire  _T_83; // @[Conditional.scala 37:30]
  wire  _GEN_6; // @[BasicBlock.scala 1045:43]
  wire  _GEN_7; // @[BasicBlock.scala 1045:43]
  wire  _GEN_8; // @[BasicBlock.scala 1066:41]
  wire [9:0] _GEN_9; // @[BasicBlock.scala 1066:41]
  wire  _GEN_10; // @[BasicBlock.scala 1066:41]
  wire  _GEN_11; // @[BasicBlock.scala 1066:41]
  wire  _GEN_12; // @[BasicBlock.scala 1066:41]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire  _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_21; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  wire  _GEN_23; // @[Conditional.scala 40:58]
  assign _T_73 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_73 ? io_predicateIn_0_bits_taskID : in_data_R_0_taskID; // @[BasicBlock.scala 998:36]
  assign _GEN_2 = _T_73 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 998:36]
  assign _GEN_3 = _T_73 ? 1'h1 : in_data_valid_R_0; // @[BasicBlock.scala 998:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 1005:34]
  assign _T_75 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_75 ? 1'h1 : output_fire_R_0; // @[BasicBlock.scala 1010:28]
  assign _GEN_5 = _T_75 ? 1'h0 : output_valid_R_0; // @[BasicBlock.scala 1010:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_75; // @[BasicBlock.scala 1027:85]
  assign _T_83 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_6 = in_data_valid_R_0 ? 1'h1 : _GEN_5; // @[BasicBlock.scala 1045:43]
  assign _GEN_7 = in_data_valid_R_0 ? 1'h1 : state; // @[BasicBlock.scala 1045:43]
  assign _GEN_8 = out_fire_mask_0 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 1066:41]
  assign _GEN_9 = out_fire_mask_0 ? 10'h0 : _GEN_1; // @[BasicBlock.scala 1066:41]
  assign _GEN_10 = out_fire_mask_0 ? 1'h0 : _GEN_3; // @[BasicBlock.scala 1066:41]
  assign _GEN_11 = out_fire_mask_0 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 1066:41]
  assign _GEN_12 = out_fire_mask_0 ? 1'h0 : state; // @[BasicBlock.scala 1066:41]
  assign _GEN_13 = state ? _GEN_8 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_14 = state ? _GEN_9 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_11 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_12 : state; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_83 ? _GEN_6 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_83 ? _GEN_7 : _GEN_17; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_83 ? _GEN_2 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_83 ? _GEN_1 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_83 ? _GEN_3 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_23 = _T_83 ? _GEN_4 : _GEN_16; // @[Conditional.scala 40:58]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 997:29]
  assign io_Out_0_valid = output_valid_R_0; // @[BasicBlock.scala 1019:21]
  assign io_Out_0_bits_taskID = output_R_taskID; // @[BasicBlock.scala 1018:20]
  assign io_Out_0_bits_control = output_R_control; // @[BasicBlock.scala 1018:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  output_R_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      in_data_R_0_taskID <= 10'h0;
    end else begin
      if (_T_83) begin
        if (_T_73) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 10'h0;
          end else begin
            if (_T_73) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_73) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_83) begin
        if (_T_73) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_73) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_73) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_83) begin
        if (_T_73) begin
          in_data_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            if (_T_73) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_73) begin
            in_data_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 10'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_R_control <= 1'h0;
    end else begin
      output_R_control <= in_data_R_0_control;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_83) begin
        if (in_data_valid_R_0) begin
          output_valid_R_0 <= 1'h1;
        end else begin
          if (_T_75) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_75) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_83) begin
        if (_T_75) begin
          output_fire_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            if (_T_75) begin
              output_fire_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_75) begin
            output_fire_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_83) begin
        if (in_data_valid_R_0) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module BasicBlockNode(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [9:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [9:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [9:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_1; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_4;
  reg  out_valid_R_2; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_5;
  reg  mask_valid_R_0; // @[HandShaking.scala 714:46]
  reg [31:0] _RAND_6;
  wire  _T_155; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 723:29]
  wire  _GEN_1; // @[HandShaking.scala 723:29]
  wire  _T_157; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 723:29]
  wire  _GEN_3; // @[HandShaking.scala 723:29]
  wire  _T_159; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 723:29]
  wire  _GEN_5; // @[HandShaking.scala 723:29]
  wire  _T_161; // @[Decoupled.scala 37:37]
  wire  _GEN_7; // @[HandShaking.scala 734:32]
  reg [9:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_7;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_8;
  reg [9:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_9;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_10;
  reg  predicate_control_R_0; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_11;
  reg  predicate_control_R_1; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_12;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_13;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_14;
  reg  state; // @[BasicBlock.scala 78:22]
  reg [31:0] _RAND_15;
  wire  _T_215; // @[Decoupled.scala 37:37]
  wire  _T_216; // @[Decoupled.scala 37:37]
  wire  _T_217; // @[BasicBlock.scala 87:91]
  wire  _T_218; // @[BasicBlock.scala 87:91]
  wire  start; // @[BasicBlock.scala 87:107]
  wire [9:0] _GEN_9; // @[BasicBlock.scala 96:36]
  wire  _GEN_10; // @[BasicBlock.scala 96:36]
  wire  _GEN_11; // @[BasicBlock.scala 96:36]
  wire  _GEN_12; // @[BasicBlock.scala 96:36]
  wire [9:0] _GEN_13; // @[BasicBlock.scala 96:36]
  wire  _GEN_14; // @[BasicBlock.scala 96:36]
  wire  _GEN_15; // @[BasicBlock.scala 96:36]
  wire  _GEN_16; // @[BasicBlock.scala 96:36]
  wire  _T_226; // @[Conditional.scala 37:30]
  wire  _GEN_17; // @[BasicBlock.scala 121:19]
  wire  _GEN_18; // @[BasicBlock.scala 121:19]
  wire  _GEN_19; // @[BasicBlock.scala 121:19]
  wire  _GEN_20; // @[BasicBlock.scala 121:19]
  wire  _GEN_21; // @[BasicBlock.scala 121:19]
  wire [2:0] _T_242; // @[HandShaking.scala 748:17]
  wire [2:0] _T_243; // @[HandShaking.scala 748:24]
  wire  _T_245; // @[HandShaking.scala 748:24]
  wire  _GEN_22; // @[BasicBlock.scala 128:26]
  wire  _GEN_23; // @[BasicBlock.scala 128:26]
  wire  _GEN_24; // @[BasicBlock.scala 128:26]
  wire  _GEN_25; // @[BasicBlock.scala 128:26]
  wire  _GEN_26; // @[BasicBlock.scala 128:26]
  wire  _GEN_28; // @[BasicBlock.scala 128:26]
  wire  _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_36; // @[Conditional.scala 40:58]
  wire  _GEN_37; // @[Conditional.scala 40:58]
  wire  _GEN_38; // @[Conditional.scala 40:58]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire  _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  assign _T_155 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_155 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 723:29]
  assign _GEN_1 = _T_155 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 723:29]
  assign _T_157 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_157 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 723:29]
  assign _GEN_3 = _T_157 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 723:29]
  assign _T_159 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_159 ? io_Out_2_ready : out_ready_R_2; // @[HandShaking.scala 723:29]
  assign _GEN_5 = _T_159 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 723:29]
  assign _T_161 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_161 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 734:32]
  assign _T_215 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _T_216 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 37:37]
  assign _T_217 = _T_215 | predicate_valid_R_0; // @[BasicBlock.scala 87:91]
  assign _T_218 = _T_216 | predicate_valid_R_1; // @[BasicBlock.scala 87:91]
  assign start = _T_217 & _T_218; // @[BasicBlock.scala 87:107]
  assign _GEN_9 = _T_215 ? io_predicateIn_0_bits_taskID : predicate_in_R_0_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_10 = _T_215 ? io_predicateIn_0_bits_control : predicate_in_R_0_control; // @[BasicBlock.scala 96:36]
  assign _GEN_11 = _T_215 ? io_predicateIn_0_bits_control : predicate_control_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_12 = _T_215 ? 1'h1 : predicate_valid_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_13 = _T_216 ? io_predicateIn_1_bits_taskID : predicate_in_R_1_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_14 = _T_216 ? io_predicateIn_1_bits_control : predicate_in_R_1_control; // @[BasicBlock.scala 96:36]
  assign _GEN_15 = _T_216 ? io_predicateIn_1_bits_control : predicate_control_R_1; // @[BasicBlock.scala 96:36]
  assign _GEN_16 = _T_216 ? 1'h1 : predicate_valid_R_1; // @[BasicBlock.scala 96:36]
  assign _T_226 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_17 = start ? 1'h1 : _GEN_1; // @[BasicBlock.scala 121:19]
  assign _GEN_18 = start ? 1'h1 : _GEN_3; // @[BasicBlock.scala 121:19]
  assign _GEN_19 = start ? 1'h1 : _GEN_5; // @[BasicBlock.scala 121:19]
  assign _GEN_20 = start ? 1'h1 : _GEN_7; // @[BasicBlock.scala 121:19]
  assign _GEN_21 = start ? 1'h1 : state; // @[BasicBlock.scala 121:19]
  assign _T_242 = {out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 748:17]
  assign _T_243 = ~ _T_242; // @[HandShaking.scala 748:24]
  assign _T_245 = _T_243 == 3'h0; // @[HandShaking.scala 748:24]
  assign _GEN_22 = _T_245 ? 1'h0 : _GEN_12; // @[BasicBlock.scala 128:26]
  assign _GEN_23 = _T_245 ? 1'h0 : _GEN_16; // @[BasicBlock.scala 128:26]
  assign _GEN_24 = _T_245 ? 1'h0 : _GEN_0; // @[BasicBlock.scala 128:26]
  assign _GEN_25 = _T_245 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 128:26]
  assign _GEN_26 = _T_245 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 128:26]
  assign _GEN_28 = _T_245 ? 1'h0 : state; // @[BasicBlock.scala 128:26]
  assign _GEN_29 = state ? _GEN_22 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_30 = state ? _GEN_23 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_31 = state ? _GEN_24 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_32 = state ? _GEN_25 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_33 = state ? _GEN_26 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_28 : state; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_226 ? _GEN_17 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_37 = _T_226 ? _GEN_18 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_38 = _T_226 ? _GEN_19 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_39 = _T_226 ? _GEN_20 : _GEN_7; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_226 ? _GEN_21 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_226 ? _GEN_12 : _GEN_29; // @[Conditional.scala 40:58]
  assign _GEN_42 = _T_226 ? _GEN_16 : _GEN_30; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_226 ? _GEN_0 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_226 ? _GEN_2 : _GEN_32; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_226 ? _GEN_4 : _GEN_33; // @[Conditional.scala 40:58]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 733:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 111:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 722:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 722:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 722:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 95:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 95:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_155) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_155) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_155) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_157) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_157) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_157) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_159) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_159) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_159) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_155) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_155) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_157) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_157) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          out_valid_R_2 <= 1'h1;
        end else begin
          if (_T_159) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_159) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          mask_valid_R_0 <= 1'h1;
        end else begin
          if (_T_161) begin
            mask_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_161) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_215) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_215) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_216) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_216) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_215) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_216) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_215) begin
          predicate_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            if (_T_215) begin
              predicate_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_215) begin
            predicate_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_216) begin
          predicate_valid_R_1 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            if (_T_216) begin
              predicate_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_216) begin
            predicate_valid_R_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module BasicBlockNode_1(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [9:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [9:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [9:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_1; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_4;
  reg  out_valid_R_2; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_5;
  reg  mask_valid_R_0; // @[HandShaking.scala 714:46]
  reg [31:0] _RAND_6;
  wire  _T_155; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 723:29]
  wire  _GEN_1; // @[HandShaking.scala 723:29]
  wire  _T_157; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 723:29]
  wire  _GEN_3; // @[HandShaking.scala 723:29]
  wire  _T_159; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 723:29]
  wire  _GEN_5; // @[HandShaking.scala 723:29]
  wire  _T_161; // @[Decoupled.scala 37:37]
  wire  _GEN_7; // @[HandShaking.scala 734:32]
  reg [9:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_7;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_8;
  reg [9:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_9;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_10;
  reg  predicate_control_R_0; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_11;
  reg  predicate_control_R_1; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_12;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_13;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_14;
  reg  state; // @[BasicBlock.scala 78:22]
  reg [31:0] _RAND_15;
  wire  _T_215; // @[Decoupled.scala 37:37]
  wire  _T_216; // @[Decoupled.scala 37:37]
  wire  _T_217; // @[BasicBlock.scala 87:91]
  wire  _T_218; // @[BasicBlock.scala 87:91]
  wire  start; // @[BasicBlock.scala 87:107]
  wire [9:0] _GEN_9; // @[BasicBlock.scala 96:36]
  wire  _GEN_10; // @[BasicBlock.scala 96:36]
  wire  _GEN_11; // @[BasicBlock.scala 96:36]
  wire  _GEN_12; // @[BasicBlock.scala 96:36]
  wire [9:0] _GEN_13; // @[BasicBlock.scala 96:36]
  wire  _GEN_14; // @[BasicBlock.scala 96:36]
  wire  _GEN_15; // @[BasicBlock.scala 96:36]
  wire  _GEN_16; // @[BasicBlock.scala 96:36]
  wire  _T_226; // @[Conditional.scala 37:30]
  wire  _GEN_17; // @[BasicBlock.scala 121:19]
  wire  _GEN_18; // @[BasicBlock.scala 121:19]
  wire  _GEN_19; // @[BasicBlock.scala 121:19]
  wire  _GEN_20; // @[BasicBlock.scala 121:19]
  wire  _GEN_21; // @[BasicBlock.scala 121:19]
  wire [2:0] _T_242; // @[HandShaking.scala 748:17]
  wire [2:0] _T_243; // @[HandShaking.scala 748:24]
  wire  _T_245; // @[HandShaking.scala 748:24]
  wire  _GEN_22; // @[BasicBlock.scala 128:26]
  wire  _GEN_23; // @[BasicBlock.scala 128:26]
  wire  _GEN_24; // @[BasicBlock.scala 128:26]
  wire  _GEN_25; // @[BasicBlock.scala 128:26]
  wire  _GEN_26; // @[BasicBlock.scala 128:26]
  wire  _GEN_28; // @[BasicBlock.scala 128:26]
  wire  _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_36; // @[Conditional.scala 40:58]
  wire  _GEN_37; // @[Conditional.scala 40:58]
  wire  _GEN_38; // @[Conditional.scala 40:58]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire  _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  assign _T_155 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_155 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 723:29]
  assign _GEN_1 = _T_155 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 723:29]
  assign _T_157 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_157 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 723:29]
  assign _GEN_3 = _T_157 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 723:29]
  assign _T_159 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_159 ? io_Out_2_ready : out_ready_R_2; // @[HandShaking.scala 723:29]
  assign _GEN_5 = _T_159 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 723:29]
  assign _T_161 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_161 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 734:32]
  assign _T_215 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _T_216 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 37:37]
  assign _T_217 = _T_215 | predicate_valid_R_0; // @[BasicBlock.scala 87:91]
  assign _T_218 = _T_216 | predicate_valid_R_1; // @[BasicBlock.scala 87:91]
  assign start = _T_217 & _T_218; // @[BasicBlock.scala 87:107]
  assign _GEN_9 = _T_215 ? io_predicateIn_0_bits_taskID : predicate_in_R_0_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_10 = _T_215 ? io_predicateIn_0_bits_control : predicate_in_R_0_control; // @[BasicBlock.scala 96:36]
  assign _GEN_11 = _T_215 ? io_predicateIn_0_bits_control : predicate_control_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_12 = _T_215 ? 1'h1 : predicate_valid_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_13 = _T_216 ? io_predicateIn_1_bits_taskID : predicate_in_R_1_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_14 = _T_216 ? io_predicateIn_1_bits_control : predicate_in_R_1_control; // @[BasicBlock.scala 96:36]
  assign _GEN_15 = _T_216 ? io_predicateIn_1_bits_control : predicate_control_R_1; // @[BasicBlock.scala 96:36]
  assign _GEN_16 = _T_216 ? 1'h1 : predicate_valid_R_1; // @[BasicBlock.scala 96:36]
  assign _T_226 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_17 = start ? 1'h1 : _GEN_1; // @[BasicBlock.scala 121:19]
  assign _GEN_18 = start ? 1'h1 : _GEN_3; // @[BasicBlock.scala 121:19]
  assign _GEN_19 = start ? 1'h1 : _GEN_5; // @[BasicBlock.scala 121:19]
  assign _GEN_20 = start ? 1'h1 : _GEN_7; // @[BasicBlock.scala 121:19]
  assign _GEN_21 = start ? 1'h1 : state; // @[BasicBlock.scala 121:19]
  assign _T_242 = {out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 748:17]
  assign _T_243 = ~ _T_242; // @[HandShaking.scala 748:24]
  assign _T_245 = _T_243 == 3'h0; // @[HandShaking.scala 748:24]
  assign _GEN_22 = _T_245 ? 1'h0 : _GEN_12; // @[BasicBlock.scala 128:26]
  assign _GEN_23 = _T_245 ? 1'h0 : _GEN_16; // @[BasicBlock.scala 128:26]
  assign _GEN_24 = _T_245 ? 1'h0 : _GEN_0; // @[BasicBlock.scala 128:26]
  assign _GEN_25 = _T_245 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 128:26]
  assign _GEN_26 = _T_245 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 128:26]
  assign _GEN_28 = _T_245 ? 1'h0 : state; // @[BasicBlock.scala 128:26]
  assign _GEN_29 = state ? _GEN_22 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_30 = state ? _GEN_23 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_31 = state ? _GEN_24 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_32 = state ? _GEN_25 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_33 = state ? _GEN_26 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_28 : state; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_226 ? _GEN_17 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_37 = _T_226 ? _GEN_18 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_38 = _T_226 ? _GEN_19 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_39 = _T_226 ? _GEN_20 : _GEN_7; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_226 ? _GEN_21 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_226 ? _GEN_12 : _GEN_29; // @[Conditional.scala 40:58]
  assign _GEN_42 = _T_226 ? _GEN_16 : _GEN_30; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_226 ? _GEN_0 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_226 ? _GEN_2 : _GEN_32; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_226 ? _GEN_4 : _GEN_33; // @[Conditional.scala 40:58]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 733:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 111:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 722:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 722:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 722:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 95:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 95:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_155) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_155) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_155) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_157) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_157) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_157) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_159) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_159) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_159) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_155) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_155) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_157) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_157) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          out_valid_R_2 <= 1'h1;
        end else begin
          if (_T_159) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_159) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          mask_valid_R_0 <= 1'h1;
        end else begin
          if (_T_161) begin
            mask_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_161) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_215) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_215) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_216) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_216) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_215) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_216) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_215) begin
          predicate_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            if (_T_215) begin
              predicate_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_215) begin
            predicate_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_226) begin
        if (_T_216) begin
          predicate_valid_R_1 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            if (_T_216) begin
              predicate_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_216) begin
            predicate_valid_R_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_226) begin
        if (start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_245) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module BasicBlockNode_2(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [9:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [9:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [9:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_6;
  reg  out_valid_R_2; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_7;
  reg  out_valid_R_3; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_8;
  reg  out_valid_R_4; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_9;
  reg  mask_valid_R_0; // @[HandShaking.scala 714:46]
  reg [31:0] _RAND_10;
  wire  _T_191; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 723:29]
  wire  _GEN_1; // @[HandShaking.scala 723:29]
  wire  _T_193; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 723:29]
  wire  _GEN_3; // @[HandShaking.scala 723:29]
  wire  _T_195; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 723:29]
  wire  _GEN_5; // @[HandShaking.scala 723:29]
  wire  _T_197; // @[Decoupled.scala 37:37]
  wire  _GEN_6; // @[HandShaking.scala 723:29]
  wire  _GEN_7; // @[HandShaking.scala 723:29]
  wire  _T_199; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[HandShaking.scala 723:29]
  wire  _GEN_9; // @[HandShaking.scala 723:29]
  wire  _T_201; // @[Decoupled.scala 37:37]
  wire  _GEN_11; // @[HandShaking.scala 734:32]
  reg [9:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_11;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_12;
  reg [9:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_13;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_14;
  reg  predicate_control_R_0; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_15;
  reg  predicate_control_R_1; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_16;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_17;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_18;
  reg  state; // @[BasicBlock.scala 78:22]
  reg [31:0] _RAND_19;
  wire  _T_255; // @[Decoupled.scala 37:37]
  wire  _T_256; // @[Decoupled.scala 37:37]
  wire  _T_257; // @[BasicBlock.scala 87:91]
  wire  _T_258; // @[BasicBlock.scala 87:91]
  wire  start; // @[BasicBlock.scala 87:107]
  wire [9:0] _GEN_13; // @[BasicBlock.scala 96:36]
  wire  _GEN_14; // @[BasicBlock.scala 96:36]
  wire  _GEN_15; // @[BasicBlock.scala 96:36]
  wire  _GEN_16; // @[BasicBlock.scala 96:36]
  wire [9:0] _GEN_17; // @[BasicBlock.scala 96:36]
  wire  _GEN_18; // @[BasicBlock.scala 96:36]
  wire  _GEN_19; // @[BasicBlock.scala 96:36]
  wire  _GEN_20; // @[BasicBlock.scala 96:36]
  wire  _T_266; // @[Conditional.scala 37:30]
  wire  _GEN_21; // @[BasicBlock.scala 121:19]
  wire  _GEN_22; // @[BasicBlock.scala 121:19]
  wire  _GEN_23; // @[BasicBlock.scala 121:19]
  wire  _GEN_24; // @[BasicBlock.scala 121:19]
  wire  _GEN_25; // @[BasicBlock.scala 121:19]
  wire  _GEN_26; // @[BasicBlock.scala 121:19]
  wire  _GEN_27; // @[BasicBlock.scala 121:19]
  wire [4:0] _T_288; // @[HandShaking.scala 748:17]
  wire [4:0] _T_289; // @[HandShaking.scala 748:24]
  wire  _T_291; // @[HandShaking.scala 748:24]
  wire  _GEN_28; // @[BasicBlock.scala 128:26]
  wire  _GEN_29; // @[BasicBlock.scala 128:26]
  wire  _GEN_30; // @[BasicBlock.scala 128:26]
  wire  _GEN_31; // @[BasicBlock.scala 128:26]
  wire  _GEN_32; // @[BasicBlock.scala 128:26]
  wire  _GEN_33; // @[BasicBlock.scala 128:26]
  wire  _GEN_34; // @[BasicBlock.scala 128:26]
  wire  _GEN_36; // @[BasicBlock.scala 128:26]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire  _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  wire  _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire  _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  wire  _GEN_56; // @[Conditional.scala 40:58]
  wire  _GEN_57; // @[Conditional.scala 40:58]
  wire  _GEN_58; // @[Conditional.scala 40:58]
  wire  _GEN_59; // @[Conditional.scala 40:58]
  assign _T_191 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_191 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 723:29]
  assign _GEN_1 = _T_191 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 723:29]
  assign _T_193 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_193 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 723:29]
  assign _GEN_3 = _T_193 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 723:29]
  assign _T_195 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_195 ? io_Out_2_ready : out_ready_R_2; // @[HandShaking.scala 723:29]
  assign _GEN_5 = _T_195 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 723:29]
  assign _T_197 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_197 ? io_Out_3_ready : out_ready_R_3; // @[HandShaking.scala 723:29]
  assign _GEN_7 = _T_197 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 723:29]
  assign _T_199 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_199 ? io_Out_4_ready : out_ready_R_4; // @[HandShaking.scala 723:29]
  assign _GEN_9 = _T_199 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 723:29]
  assign _T_201 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_201 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 734:32]
  assign _T_255 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _T_256 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 37:37]
  assign _T_257 = _T_255 | predicate_valid_R_0; // @[BasicBlock.scala 87:91]
  assign _T_258 = _T_256 | predicate_valid_R_1; // @[BasicBlock.scala 87:91]
  assign start = _T_257 & _T_258; // @[BasicBlock.scala 87:107]
  assign _GEN_13 = _T_255 ? io_predicateIn_0_bits_taskID : predicate_in_R_0_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_14 = _T_255 ? io_predicateIn_0_bits_control : predicate_in_R_0_control; // @[BasicBlock.scala 96:36]
  assign _GEN_15 = _T_255 ? io_predicateIn_0_bits_control : predicate_control_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_16 = _T_255 ? 1'h1 : predicate_valid_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_17 = _T_256 ? io_predicateIn_1_bits_taskID : predicate_in_R_1_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_18 = _T_256 ? io_predicateIn_1_bits_control : predicate_in_R_1_control; // @[BasicBlock.scala 96:36]
  assign _GEN_19 = _T_256 ? io_predicateIn_1_bits_control : predicate_control_R_1; // @[BasicBlock.scala 96:36]
  assign _GEN_20 = _T_256 ? 1'h1 : predicate_valid_R_1; // @[BasicBlock.scala 96:36]
  assign _T_266 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_21 = start ? 1'h1 : _GEN_1; // @[BasicBlock.scala 121:19]
  assign _GEN_22 = start ? 1'h1 : _GEN_3; // @[BasicBlock.scala 121:19]
  assign _GEN_23 = start ? 1'h1 : _GEN_5; // @[BasicBlock.scala 121:19]
  assign _GEN_24 = start ? 1'h1 : _GEN_7; // @[BasicBlock.scala 121:19]
  assign _GEN_25 = start ? 1'h1 : _GEN_9; // @[BasicBlock.scala 121:19]
  assign _GEN_26 = start ? 1'h1 : _GEN_11; // @[BasicBlock.scala 121:19]
  assign _GEN_27 = start ? 1'h1 : state; // @[BasicBlock.scala 121:19]
  assign _T_288 = {out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 748:17]
  assign _T_289 = ~ _T_288; // @[HandShaking.scala 748:24]
  assign _T_291 = _T_289 == 5'h0; // @[HandShaking.scala 748:24]
  assign _GEN_28 = _T_291 ? 1'h0 : _GEN_16; // @[BasicBlock.scala 128:26]
  assign _GEN_29 = _T_291 ? 1'h0 : _GEN_20; // @[BasicBlock.scala 128:26]
  assign _GEN_30 = _T_291 ? 1'h0 : _GEN_0; // @[BasicBlock.scala 128:26]
  assign _GEN_31 = _T_291 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 128:26]
  assign _GEN_32 = _T_291 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 128:26]
  assign _GEN_33 = _T_291 ? 1'h0 : _GEN_6; // @[BasicBlock.scala 128:26]
  assign _GEN_34 = _T_291 ? 1'h0 : _GEN_8; // @[BasicBlock.scala 128:26]
  assign _GEN_36 = _T_291 ? 1'h0 : state; // @[BasicBlock.scala 128:26]
  assign _GEN_37 = state ? _GEN_28 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_29 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_30 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_31 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_41 = state ? _GEN_32 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_33 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_34 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_45 = state ? _GEN_36 : state; // @[Conditional.scala 39:67]
  assign _GEN_46 = _T_266 ? _GEN_21 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_266 ? _GEN_22 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_266 ? _GEN_23 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_266 ? _GEN_24 : _GEN_7; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_266 ? _GEN_25 : _GEN_9; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_266 ? _GEN_26 : _GEN_11; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_266 ? _GEN_27 : _GEN_45; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_266 ? _GEN_16 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_266 ? _GEN_20 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_266 ? _GEN_0 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_56 = _T_266 ? _GEN_2 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_57 = _T_266 ? _GEN_4 : _GEN_41; // @[Conditional.scala 40:58]
  assign _GEN_58 = _T_266 ? _GEN_6 : _GEN_42; // @[Conditional.scala 40:58]
  assign _GEN_59 = _T_266 ? _GEN_8 : _GEN_43; // @[Conditional.scala 40:58]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 733:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 111:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 722:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 722:21]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 722:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 722:21]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 722:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 95:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 95:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_13[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  state = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_191) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_191) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_191) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_193) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_193) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_193) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_195) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_195) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_195) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_197) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_197) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_197) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_199) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_199) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_199) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_191) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_191) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_193) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_193) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          out_valid_R_2 <= 1'h1;
        end else begin
          if (_T_195) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_195) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          out_valid_R_3 <= 1'h1;
        end else begin
          if (_T_197) begin
            out_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_197) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          out_valid_R_4 <= 1'h1;
        end else begin
          if (_T_199) begin
            out_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_199) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          mask_valid_R_0 <= 1'h1;
        end else begin
          if (_T_201) begin
            mask_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_201) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_255) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_255) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_256) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_256) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_255) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_256) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_255) begin
          predicate_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            if (_T_255) begin
              predicate_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_255) begin
            predicate_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_266) begin
        if (_T_256) begin
          predicate_valid_R_1 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            if (_T_256) begin
              predicate_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_256) begin
            predicate_valid_R_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_266) begin
        if (start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_291) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module BasicBlockNode_3(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [9:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [9:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [9:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [9:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_7;
  reg  out_ready_R_8; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_8;
  reg  out_ready_R_9; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_9;
  reg  out_valid_R_0; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_10;
  reg  out_valid_R_1; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_11;
  reg  out_valid_R_2; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_12;
  reg  out_valid_R_3; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_13;
  reg  out_valid_R_4; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_14;
  reg  out_valid_R_5; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_15;
  reg  out_valid_R_6; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_16;
  reg  out_valid_R_7; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_17;
  reg  out_valid_R_8; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_18;
  reg  out_valid_R_9; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_19;
  reg  mask_valid_R_0; // @[HandShaking.scala 714:46]
  reg [31:0] _RAND_20;
  wire  _T_281; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 723:29]
  wire  _GEN_1; // @[HandShaking.scala 723:29]
  wire  _T_283; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 723:29]
  wire  _GEN_3; // @[HandShaking.scala 723:29]
  wire  _T_285; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 723:29]
  wire  _GEN_5; // @[HandShaking.scala 723:29]
  wire  _T_287; // @[Decoupled.scala 37:37]
  wire  _GEN_6; // @[HandShaking.scala 723:29]
  wire  _GEN_7; // @[HandShaking.scala 723:29]
  wire  _T_289; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[HandShaking.scala 723:29]
  wire  _GEN_9; // @[HandShaking.scala 723:29]
  wire  _T_291; // @[Decoupled.scala 37:37]
  wire  _GEN_10; // @[HandShaking.scala 723:29]
  wire  _GEN_11; // @[HandShaking.scala 723:29]
  wire  _T_293; // @[Decoupled.scala 37:37]
  wire  _GEN_12; // @[HandShaking.scala 723:29]
  wire  _GEN_13; // @[HandShaking.scala 723:29]
  wire  _T_295; // @[Decoupled.scala 37:37]
  wire  _GEN_14; // @[HandShaking.scala 723:29]
  wire  _GEN_15; // @[HandShaking.scala 723:29]
  wire  _T_297; // @[Decoupled.scala 37:37]
  wire  _GEN_16; // @[HandShaking.scala 723:29]
  wire  _GEN_17; // @[HandShaking.scala 723:29]
  wire  _T_299; // @[Decoupled.scala 37:37]
  wire  _GEN_18; // @[HandShaking.scala 723:29]
  wire  _GEN_19; // @[HandShaking.scala 723:29]
  wire  _T_301; // @[Decoupled.scala 37:37]
  wire  _GEN_21; // @[HandShaking.scala 734:32]
  reg [9:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_21;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_22;
  reg [9:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_23;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_24;
  reg  predicate_control_R_0; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_25;
  reg  predicate_control_R_1; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_26;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_27;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_28;
  reg  state; // @[BasicBlock.scala 78:22]
  reg [31:0] _RAND_29;
  wire  _T_355; // @[Decoupled.scala 37:37]
  wire  _T_356; // @[Decoupled.scala 37:37]
  wire  _T_357; // @[BasicBlock.scala 87:91]
  wire  _T_358; // @[BasicBlock.scala 87:91]
  wire  start; // @[BasicBlock.scala 87:107]
  wire [9:0] _GEN_23; // @[BasicBlock.scala 96:36]
  wire  _GEN_24; // @[BasicBlock.scala 96:36]
  wire  _GEN_25; // @[BasicBlock.scala 96:36]
  wire  _GEN_26; // @[BasicBlock.scala 96:36]
  wire [9:0] _GEN_27; // @[BasicBlock.scala 96:36]
  wire  _GEN_28; // @[BasicBlock.scala 96:36]
  wire  _GEN_29; // @[BasicBlock.scala 96:36]
  wire  _GEN_30; // @[BasicBlock.scala 96:36]
  wire  _T_366; // @[Conditional.scala 37:30]
  wire  _GEN_31; // @[BasicBlock.scala 121:19]
  wire  _GEN_32; // @[BasicBlock.scala 121:19]
  wire  _GEN_33; // @[BasicBlock.scala 121:19]
  wire  _GEN_34; // @[BasicBlock.scala 121:19]
  wire  _GEN_35; // @[BasicBlock.scala 121:19]
  wire  _GEN_36; // @[BasicBlock.scala 121:19]
  wire  _GEN_37; // @[BasicBlock.scala 121:19]
  wire  _GEN_38; // @[BasicBlock.scala 121:19]
  wire  _GEN_39; // @[BasicBlock.scala 121:19]
  wire  _GEN_40; // @[BasicBlock.scala 121:19]
  wire  _GEN_41; // @[BasicBlock.scala 121:19]
  wire  _GEN_42; // @[BasicBlock.scala 121:19]
  wire [9:0] _T_403; // @[HandShaking.scala 748:17]
  wire [9:0] _T_404; // @[HandShaking.scala 748:24]
  wire  _T_406; // @[HandShaking.scala 748:24]
  wire  _GEN_43; // @[BasicBlock.scala 128:26]
  wire  _GEN_44; // @[BasicBlock.scala 128:26]
  wire  _GEN_45; // @[BasicBlock.scala 128:26]
  wire  _GEN_46; // @[BasicBlock.scala 128:26]
  wire  _GEN_47; // @[BasicBlock.scala 128:26]
  wire  _GEN_48; // @[BasicBlock.scala 128:26]
  wire  _GEN_49; // @[BasicBlock.scala 128:26]
  wire  _GEN_50; // @[BasicBlock.scala 128:26]
  wire  _GEN_51; // @[BasicBlock.scala 128:26]
  wire  _GEN_52; // @[BasicBlock.scala 128:26]
  wire  _GEN_53; // @[BasicBlock.scala 128:26]
  wire  _GEN_54; // @[BasicBlock.scala 128:26]
  wire  _GEN_56; // @[BasicBlock.scala 128:26]
  wire  _GEN_57; // @[Conditional.scala 39:67]
  wire  _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_62; // @[Conditional.scala 39:67]
  wire  _GEN_63; // @[Conditional.scala 39:67]
  wire  _GEN_64; // @[Conditional.scala 39:67]
  wire  _GEN_65; // @[Conditional.scala 39:67]
  wire  _GEN_66; // @[Conditional.scala 39:67]
  wire  _GEN_67; // @[Conditional.scala 39:67]
  wire  _GEN_68; // @[Conditional.scala 39:67]
  wire  _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_71; // @[Conditional.scala 40:58]
  wire  _GEN_72; // @[Conditional.scala 40:58]
  wire  _GEN_73; // @[Conditional.scala 40:58]
  wire  _GEN_74; // @[Conditional.scala 40:58]
  wire  _GEN_75; // @[Conditional.scala 40:58]
  wire  _GEN_76; // @[Conditional.scala 40:58]
  wire  _GEN_77; // @[Conditional.scala 40:58]
  wire  _GEN_78; // @[Conditional.scala 40:58]
  wire  _GEN_79; // @[Conditional.scala 40:58]
  wire  _GEN_80; // @[Conditional.scala 40:58]
  wire  _GEN_81; // @[Conditional.scala 40:58]
  wire  _GEN_82; // @[Conditional.scala 40:58]
  wire  _GEN_83; // @[Conditional.scala 40:58]
  wire  _GEN_84; // @[Conditional.scala 40:58]
  wire  _GEN_85; // @[Conditional.scala 40:58]
  wire  _GEN_86; // @[Conditional.scala 40:58]
  wire  _GEN_87; // @[Conditional.scala 40:58]
  wire  _GEN_88; // @[Conditional.scala 40:58]
  wire  _GEN_89; // @[Conditional.scala 40:58]
  wire  _GEN_90; // @[Conditional.scala 40:58]
  wire  _GEN_91; // @[Conditional.scala 40:58]
  wire  _GEN_92; // @[Conditional.scala 40:58]
  wire  _GEN_93; // @[Conditional.scala 40:58]
  wire  _GEN_94; // @[Conditional.scala 40:58]
  assign _T_281 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_281 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 723:29]
  assign _GEN_1 = _T_281 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 723:29]
  assign _T_283 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_283 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 723:29]
  assign _GEN_3 = _T_283 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 723:29]
  assign _T_285 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_285 ? io_Out_2_ready : out_ready_R_2; // @[HandShaking.scala 723:29]
  assign _GEN_5 = _T_285 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 723:29]
  assign _T_287 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_287 ? io_Out_3_ready : out_ready_R_3; // @[HandShaking.scala 723:29]
  assign _GEN_7 = _T_287 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 723:29]
  assign _T_289 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_289 ? io_Out_4_ready : out_ready_R_4; // @[HandShaking.scala 723:29]
  assign _GEN_9 = _T_289 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 723:29]
  assign _T_291 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 37:37]
  assign _GEN_10 = _T_291 ? io_Out_5_ready : out_ready_R_5; // @[HandShaking.scala 723:29]
  assign _GEN_11 = _T_291 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 723:29]
  assign _T_293 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_293 ? io_Out_6_ready : out_ready_R_6; // @[HandShaking.scala 723:29]
  assign _GEN_13 = _T_293 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 723:29]
  assign _T_295 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 37:37]
  assign _GEN_14 = _T_295 ? io_Out_7_ready : out_ready_R_7; // @[HandShaking.scala 723:29]
  assign _GEN_15 = _T_295 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 723:29]
  assign _T_297 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 37:37]
  assign _GEN_16 = _T_297 ? io_Out_8_ready : out_ready_R_8; // @[HandShaking.scala 723:29]
  assign _GEN_17 = _T_297 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 723:29]
  assign _T_299 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 37:37]
  assign _GEN_18 = _T_299 ? io_Out_9_ready : out_ready_R_9; // @[HandShaking.scala 723:29]
  assign _GEN_19 = _T_299 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 723:29]
  assign _T_301 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_21 = _T_301 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 734:32]
  assign _T_355 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _T_356 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 37:37]
  assign _T_357 = _T_355 | predicate_valid_R_0; // @[BasicBlock.scala 87:91]
  assign _T_358 = _T_356 | predicate_valid_R_1; // @[BasicBlock.scala 87:91]
  assign start = _T_357 & _T_358; // @[BasicBlock.scala 87:107]
  assign _GEN_23 = _T_355 ? io_predicateIn_0_bits_taskID : predicate_in_R_0_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_24 = _T_355 ? io_predicateIn_0_bits_control : predicate_in_R_0_control; // @[BasicBlock.scala 96:36]
  assign _GEN_25 = _T_355 ? io_predicateIn_0_bits_control : predicate_control_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_26 = _T_355 ? 1'h1 : predicate_valid_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_27 = _T_356 ? io_predicateIn_1_bits_taskID : predicate_in_R_1_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_28 = _T_356 ? io_predicateIn_1_bits_control : predicate_in_R_1_control; // @[BasicBlock.scala 96:36]
  assign _GEN_29 = _T_356 ? io_predicateIn_1_bits_control : predicate_control_R_1; // @[BasicBlock.scala 96:36]
  assign _GEN_30 = _T_356 ? 1'h1 : predicate_valid_R_1; // @[BasicBlock.scala 96:36]
  assign _T_366 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_31 = start ? 1'h1 : _GEN_1; // @[BasicBlock.scala 121:19]
  assign _GEN_32 = start ? 1'h1 : _GEN_3; // @[BasicBlock.scala 121:19]
  assign _GEN_33 = start ? 1'h1 : _GEN_5; // @[BasicBlock.scala 121:19]
  assign _GEN_34 = start ? 1'h1 : _GEN_7; // @[BasicBlock.scala 121:19]
  assign _GEN_35 = start ? 1'h1 : _GEN_9; // @[BasicBlock.scala 121:19]
  assign _GEN_36 = start ? 1'h1 : _GEN_11; // @[BasicBlock.scala 121:19]
  assign _GEN_37 = start ? 1'h1 : _GEN_13; // @[BasicBlock.scala 121:19]
  assign _GEN_38 = start ? 1'h1 : _GEN_15; // @[BasicBlock.scala 121:19]
  assign _GEN_39 = start ? 1'h1 : _GEN_17; // @[BasicBlock.scala 121:19]
  assign _GEN_40 = start ? 1'h1 : _GEN_19; // @[BasicBlock.scala 121:19]
  assign _GEN_41 = start ? 1'h1 : _GEN_21; // @[BasicBlock.scala 121:19]
  assign _GEN_42 = start ? 1'h1 : state; // @[BasicBlock.scala 121:19]
  assign _T_403 = {out_ready_R_9,out_ready_R_8,out_ready_R_7,out_ready_R_6,out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 748:17]
  assign _T_404 = ~ _T_403; // @[HandShaking.scala 748:24]
  assign _T_406 = _T_404 == 10'h0; // @[HandShaking.scala 748:24]
  assign _GEN_43 = _T_406 ? 1'h0 : _GEN_26; // @[BasicBlock.scala 128:26]
  assign _GEN_44 = _T_406 ? 1'h0 : _GEN_30; // @[BasicBlock.scala 128:26]
  assign _GEN_45 = _T_406 ? 1'h0 : _GEN_0; // @[BasicBlock.scala 128:26]
  assign _GEN_46 = _T_406 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 128:26]
  assign _GEN_47 = _T_406 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 128:26]
  assign _GEN_48 = _T_406 ? 1'h0 : _GEN_6; // @[BasicBlock.scala 128:26]
  assign _GEN_49 = _T_406 ? 1'h0 : _GEN_8; // @[BasicBlock.scala 128:26]
  assign _GEN_50 = _T_406 ? 1'h0 : _GEN_10; // @[BasicBlock.scala 128:26]
  assign _GEN_51 = _T_406 ? 1'h0 : _GEN_12; // @[BasicBlock.scala 128:26]
  assign _GEN_52 = _T_406 ? 1'h0 : _GEN_14; // @[BasicBlock.scala 128:26]
  assign _GEN_53 = _T_406 ? 1'h0 : _GEN_16; // @[BasicBlock.scala 128:26]
  assign _GEN_54 = _T_406 ? 1'h0 : _GEN_18; // @[BasicBlock.scala 128:26]
  assign _GEN_56 = _T_406 ? 1'h0 : state; // @[BasicBlock.scala 128:26]
  assign _GEN_57 = state ? _GEN_43 : _GEN_26; // @[Conditional.scala 39:67]
  assign _GEN_58 = state ? _GEN_44 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_59 = state ? _GEN_45 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_60 = state ? _GEN_46 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_61 = state ? _GEN_47 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_62 = state ? _GEN_48 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_63 = state ? _GEN_49 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_64 = state ? _GEN_50 : _GEN_10; // @[Conditional.scala 39:67]
  assign _GEN_65 = state ? _GEN_51 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_66 = state ? _GEN_52 : _GEN_14; // @[Conditional.scala 39:67]
  assign _GEN_67 = state ? _GEN_53 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_68 = state ? _GEN_54 : _GEN_18; // @[Conditional.scala 39:67]
  assign _GEN_70 = state ? _GEN_56 : state; // @[Conditional.scala 39:67]
  assign _GEN_71 = _T_366 ? _GEN_31 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_72 = _T_366 ? _GEN_32 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_73 = _T_366 ? _GEN_33 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_74 = _T_366 ? _GEN_34 : _GEN_7; // @[Conditional.scala 40:58]
  assign _GEN_75 = _T_366 ? _GEN_35 : _GEN_9; // @[Conditional.scala 40:58]
  assign _GEN_76 = _T_366 ? _GEN_36 : _GEN_11; // @[Conditional.scala 40:58]
  assign _GEN_77 = _T_366 ? _GEN_37 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_78 = _T_366 ? _GEN_38 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_79 = _T_366 ? _GEN_39 : _GEN_17; // @[Conditional.scala 40:58]
  assign _GEN_80 = _T_366 ? _GEN_40 : _GEN_19; // @[Conditional.scala 40:58]
  assign _GEN_81 = _T_366 ? _GEN_41 : _GEN_21; // @[Conditional.scala 40:58]
  assign _GEN_82 = _T_366 ? _GEN_42 : _GEN_70; // @[Conditional.scala 40:58]
  assign _GEN_83 = _T_366 ? _GEN_26 : _GEN_57; // @[Conditional.scala 40:58]
  assign _GEN_84 = _T_366 ? _GEN_30 : _GEN_58; // @[Conditional.scala 40:58]
  assign _GEN_85 = _T_366 ? _GEN_0 : _GEN_59; // @[Conditional.scala 40:58]
  assign _GEN_86 = _T_366 ? _GEN_2 : _GEN_60; // @[Conditional.scala 40:58]
  assign _GEN_87 = _T_366 ? _GEN_4 : _GEN_61; // @[Conditional.scala 40:58]
  assign _GEN_88 = _T_366 ? _GEN_6 : _GEN_62; // @[Conditional.scala 40:58]
  assign _GEN_89 = _T_366 ? _GEN_8 : _GEN_63; // @[Conditional.scala 40:58]
  assign _GEN_90 = _T_366 ? _GEN_10 : _GEN_64; // @[Conditional.scala 40:58]
  assign _GEN_91 = _T_366 ? _GEN_12 : _GEN_65; // @[Conditional.scala 40:58]
  assign _GEN_92 = _T_366 ? _GEN_14 : _GEN_66; // @[Conditional.scala 40:58]
  assign _GEN_93 = _T_366 ? _GEN_16 : _GEN_67; // @[Conditional.scala 40:58]
  assign _GEN_94 = _T_366 ? _GEN_18 : _GEN_68; // @[Conditional.scala 40:58]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 733:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 111:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 722:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 722:21]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 722:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 722:21]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 722:21]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 722:21]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 722:21]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 722:21]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 722:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_8_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 722:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_9_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 95:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 95:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_21[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_23[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  state = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_281) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_281) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_281) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_283) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_283) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_283) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_285) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_285) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_285) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_287) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_287) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_287) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_289) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_289) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_289) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_291) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_291) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_291) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_293) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_293) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_293) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_295) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_295) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_295) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_297) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_297) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_297) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_299) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_299) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_299) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_281) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_281) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_283) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_283) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_2 <= 1'h1;
        end else begin
          if (_T_285) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_285) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_3 <= 1'h1;
        end else begin
          if (_T_287) begin
            out_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_287) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_4 <= 1'h1;
        end else begin
          if (_T_289) begin
            out_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_289) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_5 <= 1'h1;
        end else begin
          if (_T_291) begin
            out_valid_R_5 <= 1'h0;
          end
        end
      end else begin
        if (_T_291) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_6 <= 1'h1;
        end else begin
          if (_T_293) begin
            out_valid_R_6 <= 1'h0;
          end
        end
      end else begin
        if (_T_293) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_7 <= 1'h1;
        end else begin
          if (_T_295) begin
            out_valid_R_7 <= 1'h0;
          end
        end
      end else begin
        if (_T_295) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_8 <= 1'h1;
        end else begin
          if (_T_297) begin
            out_valid_R_8 <= 1'h0;
          end
        end
      end else begin
        if (_T_297) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          out_valid_R_9 <= 1'h1;
        end else begin
          if (_T_299) begin
            out_valid_R_9 <= 1'h0;
          end
        end
      end else begin
        if (_T_299) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          mask_valid_R_0 <= 1'h1;
        end else begin
          if (_T_301) begin
            mask_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_301) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_355) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_355) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_356) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_356) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_355) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_356) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_355) begin
          predicate_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            if (_T_355) begin
              predicate_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_355) begin
            predicate_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_366) begin
        if (_T_356) begin
          predicate_valid_R_1 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            if (_T_356) begin
              predicate_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_356) begin
            predicate_valid_R_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_366) begin
        if (start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_406) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module BasicBlockNode_4(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [9:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [9:0] io_Out_2_bits_taskID,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [9:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [9:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [9:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output       io_Out_9_bits_control,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output       io_Out_10_bits_control,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output       io_Out_11_bits_control,
  input        io_Out_12_ready,
  output       io_Out_12_valid,
  output [9:0] io_Out_12_bits_taskID,
  output       io_Out_12_bits_control,
  input        io_Out_13_ready,
  output       io_Out_13_valid,
  output [9:0] io_Out_13_bits_taskID,
  output       io_Out_13_bits_control,
  input        io_Out_14_ready,
  output       io_Out_14_valid,
  output [9:0] io_Out_14_bits_taskID,
  output       io_Out_14_bits_control,
  input        io_Out_15_ready,
  output       io_Out_15_valid,
  output [9:0] io_Out_15_bits_taskID,
  output       io_Out_15_bits_control,
  input        io_Out_16_ready,
  output       io_Out_16_valid,
  output [9:0] io_Out_16_bits_taskID,
  output       io_Out_16_bits_control,
  input        io_Out_17_ready,
  output       io_Out_17_valid,
  output [9:0] io_Out_17_bits_taskID,
  output       io_Out_17_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [9:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_7;
  reg  out_ready_R_8; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_8;
  reg  out_ready_R_9; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_9;
  reg  out_ready_R_10; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_10;
  reg  out_ready_R_11; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_11;
  reg  out_ready_R_12; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_12;
  reg  out_ready_R_13; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_13;
  reg  out_ready_R_14; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_14;
  reg  out_ready_R_15; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_15;
  reg  out_ready_R_16; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_16;
  reg  out_ready_R_17; // @[HandShaking.scala 709:28]
  reg [31:0] _RAND_17;
  reg  out_valid_R_0; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_18;
  reg  out_valid_R_1; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_19;
  reg  out_valid_R_2; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_20;
  reg  out_valid_R_3; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_21;
  reg  out_valid_R_4; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_22;
  reg  out_valid_R_5; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_23;
  reg  out_valid_R_6; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_24;
  reg  out_valid_R_7; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_25;
  reg  out_valid_R_8; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_26;
  reg  out_valid_R_9; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_27;
  reg  out_valid_R_10; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_28;
  reg  out_valid_R_11; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_29;
  reg  out_valid_R_12; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_30;
  reg  out_valid_R_13; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_31;
  reg  out_valid_R_14; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_32;
  reg  out_valid_R_15; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_33;
  reg  out_valid_R_16; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_34;
  reg  out_valid_R_17; // @[HandShaking.scala 710:28]
  reg [31:0] _RAND_35;
  reg  mask_valid_R_0; // @[HandShaking.scala 714:46]
  reg [31:0] _RAND_36;
  wire  _T_425; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 723:29]
  wire  _GEN_1; // @[HandShaking.scala 723:29]
  wire  _T_427; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 723:29]
  wire  _GEN_3; // @[HandShaking.scala 723:29]
  wire  _T_429; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 723:29]
  wire  _GEN_5; // @[HandShaking.scala 723:29]
  wire  _T_431; // @[Decoupled.scala 37:37]
  wire  _GEN_6; // @[HandShaking.scala 723:29]
  wire  _GEN_7; // @[HandShaking.scala 723:29]
  wire  _T_433; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[HandShaking.scala 723:29]
  wire  _GEN_9; // @[HandShaking.scala 723:29]
  wire  _T_435; // @[Decoupled.scala 37:37]
  wire  _GEN_10; // @[HandShaking.scala 723:29]
  wire  _GEN_11; // @[HandShaking.scala 723:29]
  wire  _T_437; // @[Decoupled.scala 37:37]
  wire  _GEN_12; // @[HandShaking.scala 723:29]
  wire  _GEN_13; // @[HandShaking.scala 723:29]
  wire  _T_439; // @[Decoupled.scala 37:37]
  wire  _GEN_14; // @[HandShaking.scala 723:29]
  wire  _GEN_15; // @[HandShaking.scala 723:29]
  wire  _T_441; // @[Decoupled.scala 37:37]
  wire  _GEN_16; // @[HandShaking.scala 723:29]
  wire  _GEN_17; // @[HandShaking.scala 723:29]
  wire  _T_443; // @[Decoupled.scala 37:37]
  wire  _GEN_18; // @[HandShaking.scala 723:29]
  wire  _GEN_19; // @[HandShaking.scala 723:29]
  wire  _T_445; // @[Decoupled.scala 37:37]
  wire  _GEN_20; // @[HandShaking.scala 723:29]
  wire  _GEN_21; // @[HandShaking.scala 723:29]
  wire  _T_447; // @[Decoupled.scala 37:37]
  wire  _GEN_22; // @[HandShaking.scala 723:29]
  wire  _GEN_23; // @[HandShaking.scala 723:29]
  wire  _T_449; // @[Decoupled.scala 37:37]
  wire  _GEN_24; // @[HandShaking.scala 723:29]
  wire  _GEN_25; // @[HandShaking.scala 723:29]
  wire  _T_451; // @[Decoupled.scala 37:37]
  wire  _GEN_26; // @[HandShaking.scala 723:29]
  wire  _GEN_27; // @[HandShaking.scala 723:29]
  wire  _T_453; // @[Decoupled.scala 37:37]
  wire  _GEN_28; // @[HandShaking.scala 723:29]
  wire  _GEN_29; // @[HandShaking.scala 723:29]
  wire  _T_455; // @[Decoupled.scala 37:37]
  wire  _GEN_30; // @[HandShaking.scala 723:29]
  wire  _GEN_31; // @[HandShaking.scala 723:29]
  wire  _T_457; // @[Decoupled.scala 37:37]
  wire  _GEN_32; // @[HandShaking.scala 723:29]
  wire  _GEN_33; // @[HandShaking.scala 723:29]
  wire  _T_459; // @[Decoupled.scala 37:37]
  wire  _GEN_34; // @[HandShaking.scala 723:29]
  wire  _GEN_35; // @[HandShaking.scala 723:29]
  wire  _T_461; // @[Decoupled.scala 37:37]
  wire  _GEN_37; // @[HandShaking.scala 734:32]
  reg [9:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_37;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_38;
  reg [9:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_39;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 73:51]
  reg [31:0] _RAND_40;
  reg  predicate_control_R_0; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_41;
  reg  predicate_control_R_1; // @[BasicBlock.scala 74:36]
  reg [31:0] _RAND_42;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_43;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 75:54]
  reg [31:0] _RAND_44;
  reg  state; // @[BasicBlock.scala 78:22]
  reg [31:0] _RAND_45;
  wire  _T_515; // @[Decoupled.scala 37:37]
  wire  _T_516; // @[Decoupled.scala 37:37]
  wire  _T_517; // @[BasicBlock.scala 87:91]
  wire  _T_518; // @[BasicBlock.scala 87:91]
  wire  start; // @[BasicBlock.scala 87:107]
  wire [9:0] _GEN_39; // @[BasicBlock.scala 96:36]
  wire  _GEN_40; // @[BasicBlock.scala 96:36]
  wire  _GEN_41; // @[BasicBlock.scala 96:36]
  wire  _GEN_42; // @[BasicBlock.scala 96:36]
  wire [9:0] _GEN_43; // @[BasicBlock.scala 96:36]
  wire  _GEN_44; // @[BasicBlock.scala 96:36]
  wire  _GEN_45; // @[BasicBlock.scala 96:36]
  wire  _GEN_46; // @[BasicBlock.scala 96:36]
  wire  _T_526; // @[Conditional.scala 37:30]
  wire  _GEN_47; // @[BasicBlock.scala 121:19]
  wire  _GEN_48; // @[BasicBlock.scala 121:19]
  wire  _GEN_49; // @[BasicBlock.scala 121:19]
  wire  _GEN_50; // @[BasicBlock.scala 121:19]
  wire  _GEN_51; // @[BasicBlock.scala 121:19]
  wire  _GEN_52; // @[BasicBlock.scala 121:19]
  wire  _GEN_53; // @[BasicBlock.scala 121:19]
  wire  _GEN_54; // @[BasicBlock.scala 121:19]
  wire  _GEN_55; // @[BasicBlock.scala 121:19]
  wire  _GEN_56; // @[BasicBlock.scala 121:19]
  wire  _GEN_57; // @[BasicBlock.scala 121:19]
  wire  _GEN_58; // @[BasicBlock.scala 121:19]
  wire  _GEN_59; // @[BasicBlock.scala 121:19]
  wire  _GEN_60; // @[BasicBlock.scala 121:19]
  wire  _GEN_61; // @[BasicBlock.scala 121:19]
  wire  _GEN_62; // @[BasicBlock.scala 121:19]
  wire  _GEN_63; // @[BasicBlock.scala 121:19]
  wire  _GEN_64; // @[BasicBlock.scala 121:19]
  wire  _GEN_65; // @[BasicBlock.scala 121:19]
  wire  _GEN_66; // @[BasicBlock.scala 121:19]
  wire [8:0] _T_578; // @[HandShaking.scala 748:17]
  wire [17:0] _T_587; // @[HandShaking.scala 748:17]
  wire [17:0] _T_588; // @[HandShaking.scala 748:24]
  wire  _T_590; // @[HandShaking.scala 748:24]
  wire  _GEN_67; // @[BasicBlock.scala 128:26]
  wire  _GEN_68; // @[BasicBlock.scala 128:26]
  wire  _GEN_69; // @[BasicBlock.scala 128:26]
  wire  _GEN_70; // @[BasicBlock.scala 128:26]
  wire  _GEN_71; // @[BasicBlock.scala 128:26]
  wire  _GEN_72; // @[BasicBlock.scala 128:26]
  wire  _GEN_73; // @[BasicBlock.scala 128:26]
  wire  _GEN_74; // @[BasicBlock.scala 128:26]
  wire  _GEN_75; // @[BasicBlock.scala 128:26]
  wire  _GEN_76; // @[BasicBlock.scala 128:26]
  wire  _GEN_77; // @[BasicBlock.scala 128:26]
  wire  _GEN_78; // @[BasicBlock.scala 128:26]
  wire  _GEN_79; // @[BasicBlock.scala 128:26]
  wire  _GEN_80; // @[BasicBlock.scala 128:26]
  wire  _GEN_81; // @[BasicBlock.scala 128:26]
  wire  _GEN_82; // @[BasicBlock.scala 128:26]
  wire  _GEN_83; // @[BasicBlock.scala 128:26]
  wire  _GEN_84; // @[BasicBlock.scala 128:26]
  wire  _GEN_85; // @[BasicBlock.scala 128:26]
  wire  _GEN_86; // @[BasicBlock.scala 128:26]
  wire  _GEN_88; // @[BasicBlock.scala 128:26]
  wire  _GEN_89; // @[Conditional.scala 39:67]
  wire  _GEN_90; // @[Conditional.scala 39:67]
  wire  _GEN_91; // @[Conditional.scala 39:67]
  wire  _GEN_92; // @[Conditional.scala 39:67]
  wire  _GEN_93; // @[Conditional.scala 39:67]
  wire  _GEN_94; // @[Conditional.scala 39:67]
  wire  _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_96; // @[Conditional.scala 39:67]
  wire  _GEN_97; // @[Conditional.scala 39:67]
  wire  _GEN_98; // @[Conditional.scala 39:67]
  wire  _GEN_99; // @[Conditional.scala 39:67]
  wire  _GEN_100; // @[Conditional.scala 39:67]
  wire  _GEN_101; // @[Conditional.scala 39:67]
  wire  _GEN_102; // @[Conditional.scala 39:67]
  wire  _GEN_103; // @[Conditional.scala 39:67]
  wire  _GEN_104; // @[Conditional.scala 39:67]
  wire  _GEN_105; // @[Conditional.scala 39:67]
  wire  _GEN_106; // @[Conditional.scala 39:67]
  wire  _GEN_107; // @[Conditional.scala 39:67]
  wire  _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_110; // @[Conditional.scala 39:67]
  wire  _GEN_111; // @[Conditional.scala 40:58]
  wire  _GEN_112; // @[Conditional.scala 40:58]
  wire  _GEN_113; // @[Conditional.scala 40:58]
  wire  _GEN_114; // @[Conditional.scala 40:58]
  wire  _GEN_115; // @[Conditional.scala 40:58]
  wire  _GEN_116; // @[Conditional.scala 40:58]
  wire  _GEN_117; // @[Conditional.scala 40:58]
  wire  _GEN_118; // @[Conditional.scala 40:58]
  wire  _GEN_119; // @[Conditional.scala 40:58]
  wire  _GEN_120; // @[Conditional.scala 40:58]
  wire  _GEN_121; // @[Conditional.scala 40:58]
  wire  _GEN_122; // @[Conditional.scala 40:58]
  wire  _GEN_123; // @[Conditional.scala 40:58]
  wire  _GEN_124; // @[Conditional.scala 40:58]
  wire  _GEN_125; // @[Conditional.scala 40:58]
  wire  _GEN_126; // @[Conditional.scala 40:58]
  wire  _GEN_127; // @[Conditional.scala 40:58]
  wire  _GEN_128; // @[Conditional.scala 40:58]
  wire  _GEN_129; // @[Conditional.scala 40:58]
  wire  _GEN_130; // @[Conditional.scala 40:58]
  wire  _GEN_131; // @[Conditional.scala 40:58]
  wire  _GEN_132; // @[Conditional.scala 40:58]
  wire  _GEN_133; // @[Conditional.scala 40:58]
  wire  _GEN_134; // @[Conditional.scala 40:58]
  wire  _GEN_135; // @[Conditional.scala 40:58]
  wire  _GEN_136; // @[Conditional.scala 40:58]
  wire  _GEN_137; // @[Conditional.scala 40:58]
  wire  _GEN_138; // @[Conditional.scala 40:58]
  wire  _GEN_139; // @[Conditional.scala 40:58]
  wire  _GEN_140; // @[Conditional.scala 40:58]
  wire  _GEN_141; // @[Conditional.scala 40:58]
  wire  _GEN_142; // @[Conditional.scala 40:58]
  wire  _GEN_143; // @[Conditional.scala 40:58]
  wire  _GEN_144; // @[Conditional.scala 40:58]
  wire  _GEN_145; // @[Conditional.scala 40:58]
  wire  _GEN_146; // @[Conditional.scala 40:58]
  wire  _GEN_147; // @[Conditional.scala 40:58]
  wire  _GEN_148; // @[Conditional.scala 40:58]
  wire  _GEN_149; // @[Conditional.scala 40:58]
  wire  _GEN_150; // @[Conditional.scala 40:58]
  assign _T_425 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_425 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 723:29]
  assign _GEN_1 = _T_425 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 723:29]
  assign _T_427 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_427 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 723:29]
  assign _GEN_3 = _T_427 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 723:29]
  assign _T_429 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_429 ? io_Out_2_ready : out_ready_R_2; // @[HandShaking.scala 723:29]
  assign _GEN_5 = _T_429 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 723:29]
  assign _T_431 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_431 ? io_Out_3_ready : out_ready_R_3; // @[HandShaking.scala 723:29]
  assign _GEN_7 = _T_431 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 723:29]
  assign _T_433 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_433 ? io_Out_4_ready : out_ready_R_4; // @[HandShaking.scala 723:29]
  assign _GEN_9 = _T_433 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 723:29]
  assign _T_435 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 37:37]
  assign _GEN_10 = _T_435 ? io_Out_5_ready : out_ready_R_5; // @[HandShaking.scala 723:29]
  assign _GEN_11 = _T_435 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 723:29]
  assign _T_437 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_437 ? io_Out_6_ready : out_ready_R_6; // @[HandShaking.scala 723:29]
  assign _GEN_13 = _T_437 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 723:29]
  assign _T_439 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 37:37]
  assign _GEN_14 = _T_439 ? io_Out_7_ready : out_ready_R_7; // @[HandShaking.scala 723:29]
  assign _GEN_15 = _T_439 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 723:29]
  assign _T_441 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 37:37]
  assign _GEN_16 = _T_441 ? io_Out_8_ready : out_ready_R_8; // @[HandShaking.scala 723:29]
  assign _GEN_17 = _T_441 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 723:29]
  assign _T_443 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 37:37]
  assign _GEN_18 = _T_443 ? io_Out_9_ready : out_ready_R_9; // @[HandShaking.scala 723:29]
  assign _GEN_19 = _T_443 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 723:29]
  assign _T_445 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 37:37]
  assign _GEN_20 = _T_445 ? io_Out_10_ready : out_ready_R_10; // @[HandShaking.scala 723:29]
  assign _GEN_21 = _T_445 ? 1'h0 : out_valid_R_10; // @[HandShaking.scala 723:29]
  assign _T_447 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 37:37]
  assign _GEN_22 = _T_447 ? io_Out_11_ready : out_ready_R_11; // @[HandShaking.scala 723:29]
  assign _GEN_23 = _T_447 ? 1'h0 : out_valid_R_11; // @[HandShaking.scala 723:29]
  assign _T_449 = io_Out_12_ready & io_Out_12_valid; // @[Decoupled.scala 37:37]
  assign _GEN_24 = _T_449 ? io_Out_12_ready : out_ready_R_12; // @[HandShaking.scala 723:29]
  assign _GEN_25 = _T_449 ? 1'h0 : out_valid_R_12; // @[HandShaking.scala 723:29]
  assign _T_451 = io_Out_13_ready & io_Out_13_valid; // @[Decoupled.scala 37:37]
  assign _GEN_26 = _T_451 ? io_Out_13_ready : out_ready_R_13; // @[HandShaking.scala 723:29]
  assign _GEN_27 = _T_451 ? 1'h0 : out_valid_R_13; // @[HandShaking.scala 723:29]
  assign _T_453 = io_Out_14_ready & io_Out_14_valid; // @[Decoupled.scala 37:37]
  assign _GEN_28 = _T_453 ? io_Out_14_ready : out_ready_R_14; // @[HandShaking.scala 723:29]
  assign _GEN_29 = _T_453 ? 1'h0 : out_valid_R_14; // @[HandShaking.scala 723:29]
  assign _T_455 = io_Out_15_ready & io_Out_15_valid; // @[Decoupled.scala 37:37]
  assign _GEN_30 = _T_455 ? io_Out_15_ready : out_ready_R_15; // @[HandShaking.scala 723:29]
  assign _GEN_31 = _T_455 ? 1'h0 : out_valid_R_15; // @[HandShaking.scala 723:29]
  assign _T_457 = io_Out_16_ready & io_Out_16_valid; // @[Decoupled.scala 37:37]
  assign _GEN_32 = _T_457 ? io_Out_16_ready : out_ready_R_16; // @[HandShaking.scala 723:29]
  assign _GEN_33 = _T_457 ? 1'h0 : out_valid_R_16; // @[HandShaking.scala 723:29]
  assign _T_459 = io_Out_17_ready & io_Out_17_valid; // @[Decoupled.scala 37:37]
  assign _GEN_34 = _T_459 ? io_Out_17_ready : out_ready_R_17; // @[HandShaking.scala 723:29]
  assign _GEN_35 = _T_459 ? 1'h0 : out_valid_R_17; // @[HandShaking.scala 723:29]
  assign _T_461 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_37 = _T_461 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 734:32]
  assign _T_515 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _T_516 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 37:37]
  assign _T_517 = _T_515 | predicate_valid_R_0; // @[BasicBlock.scala 87:91]
  assign _T_518 = _T_516 | predicate_valid_R_1; // @[BasicBlock.scala 87:91]
  assign start = _T_517 & _T_518; // @[BasicBlock.scala 87:107]
  assign _GEN_39 = _T_515 ? io_predicateIn_0_bits_taskID : predicate_in_R_0_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_40 = _T_515 ? io_predicateIn_0_bits_control : predicate_in_R_0_control; // @[BasicBlock.scala 96:36]
  assign _GEN_41 = _T_515 ? io_predicateIn_0_bits_control : predicate_control_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_42 = _T_515 ? 1'h1 : predicate_valid_R_0; // @[BasicBlock.scala 96:36]
  assign _GEN_43 = _T_516 ? io_predicateIn_1_bits_taskID : predicate_in_R_1_taskID; // @[BasicBlock.scala 96:36]
  assign _GEN_44 = _T_516 ? io_predicateIn_1_bits_control : predicate_in_R_1_control; // @[BasicBlock.scala 96:36]
  assign _GEN_45 = _T_516 ? io_predicateIn_1_bits_control : predicate_control_R_1; // @[BasicBlock.scala 96:36]
  assign _GEN_46 = _T_516 ? 1'h1 : predicate_valid_R_1; // @[BasicBlock.scala 96:36]
  assign _T_526 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_47 = start ? 1'h1 : _GEN_1; // @[BasicBlock.scala 121:19]
  assign _GEN_48 = start ? 1'h1 : _GEN_3; // @[BasicBlock.scala 121:19]
  assign _GEN_49 = start ? 1'h1 : _GEN_5; // @[BasicBlock.scala 121:19]
  assign _GEN_50 = start ? 1'h1 : _GEN_7; // @[BasicBlock.scala 121:19]
  assign _GEN_51 = start ? 1'h1 : _GEN_9; // @[BasicBlock.scala 121:19]
  assign _GEN_52 = start ? 1'h1 : _GEN_11; // @[BasicBlock.scala 121:19]
  assign _GEN_53 = start ? 1'h1 : _GEN_13; // @[BasicBlock.scala 121:19]
  assign _GEN_54 = start ? 1'h1 : _GEN_15; // @[BasicBlock.scala 121:19]
  assign _GEN_55 = start ? 1'h1 : _GEN_17; // @[BasicBlock.scala 121:19]
  assign _GEN_56 = start ? 1'h1 : _GEN_19; // @[BasicBlock.scala 121:19]
  assign _GEN_57 = start ? 1'h1 : _GEN_21; // @[BasicBlock.scala 121:19]
  assign _GEN_58 = start ? 1'h1 : _GEN_23; // @[BasicBlock.scala 121:19]
  assign _GEN_59 = start ? 1'h1 : _GEN_25; // @[BasicBlock.scala 121:19]
  assign _GEN_60 = start ? 1'h1 : _GEN_27; // @[BasicBlock.scala 121:19]
  assign _GEN_61 = start ? 1'h1 : _GEN_29; // @[BasicBlock.scala 121:19]
  assign _GEN_62 = start ? 1'h1 : _GEN_31; // @[BasicBlock.scala 121:19]
  assign _GEN_63 = start ? 1'h1 : _GEN_33; // @[BasicBlock.scala 121:19]
  assign _GEN_64 = start ? 1'h1 : _GEN_35; // @[BasicBlock.scala 121:19]
  assign _GEN_65 = start ? 1'h1 : _GEN_37; // @[BasicBlock.scala 121:19]
  assign _GEN_66 = start ? 1'h1 : state; // @[BasicBlock.scala 121:19]
  assign _T_578 = {out_ready_R_8,out_ready_R_7,out_ready_R_6,out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 748:17]
  assign _T_587 = {out_ready_R_17,out_ready_R_16,out_ready_R_15,out_ready_R_14,out_ready_R_13,out_ready_R_12,out_ready_R_11,out_ready_R_10,out_ready_R_9,_T_578}; // @[HandShaking.scala 748:17]
  assign _T_588 = ~ _T_587; // @[HandShaking.scala 748:24]
  assign _T_590 = _T_588 == 18'h0; // @[HandShaking.scala 748:24]
  assign _GEN_67 = _T_590 ? 1'h0 : _GEN_42; // @[BasicBlock.scala 128:26]
  assign _GEN_68 = _T_590 ? 1'h0 : _GEN_46; // @[BasicBlock.scala 128:26]
  assign _GEN_69 = _T_590 ? 1'h0 : _GEN_0; // @[BasicBlock.scala 128:26]
  assign _GEN_70 = _T_590 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 128:26]
  assign _GEN_71 = _T_590 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 128:26]
  assign _GEN_72 = _T_590 ? 1'h0 : _GEN_6; // @[BasicBlock.scala 128:26]
  assign _GEN_73 = _T_590 ? 1'h0 : _GEN_8; // @[BasicBlock.scala 128:26]
  assign _GEN_74 = _T_590 ? 1'h0 : _GEN_10; // @[BasicBlock.scala 128:26]
  assign _GEN_75 = _T_590 ? 1'h0 : _GEN_12; // @[BasicBlock.scala 128:26]
  assign _GEN_76 = _T_590 ? 1'h0 : _GEN_14; // @[BasicBlock.scala 128:26]
  assign _GEN_77 = _T_590 ? 1'h0 : _GEN_16; // @[BasicBlock.scala 128:26]
  assign _GEN_78 = _T_590 ? 1'h0 : _GEN_18; // @[BasicBlock.scala 128:26]
  assign _GEN_79 = _T_590 ? 1'h0 : _GEN_20; // @[BasicBlock.scala 128:26]
  assign _GEN_80 = _T_590 ? 1'h0 : _GEN_22; // @[BasicBlock.scala 128:26]
  assign _GEN_81 = _T_590 ? 1'h0 : _GEN_24; // @[BasicBlock.scala 128:26]
  assign _GEN_82 = _T_590 ? 1'h0 : _GEN_26; // @[BasicBlock.scala 128:26]
  assign _GEN_83 = _T_590 ? 1'h0 : _GEN_28; // @[BasicBlock.scala 128:26]
  assign _GEN_84 = _T_590 ? 1'h0 : _GEN_30; // @[BasicBlock.scala 128:26]
  assign _GEN_85 = _T_590 ? 1'h0 : _GEN_32; // @[BasicBlock.scala 128:26]
  assign _GEN_86 = _T_590 ? 1'h0 : _GEN_34; // @[BasicBlock.scala 128:26]
  assign _GEN_88 = _T_590 ? 1'h0 : state; // @[BasicBlock.scala 128:26]
  assign _GEN_89 = state ? _GEN_67 : _GEN_42; // @[Conditional.scala 39:67]
  assign _GEN_90 = state ? _GEN_68 : _GEN_46; // @[Conditional.scala 39:67]
  assign _GEN_91 = state ? _GEN_69 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_92 = state ? _GEN_70 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_93 = state ? _GEN_71 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_94 = state ? _GEN_72 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_95 = state ? _GEN_73 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_96 = state ? _GEN_74 : _GEN_10; // @[Conditional.scala 39:67]
  assign _GEN_97 = state ? _GEN_75 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_98 = state ? _GEN_76 : _GEN_14; // @[Conditional.scala 39:67]
  assign _GEN_99 = state ? _GEN_77 : _GEN_16; // @[Conditional.scala 39:67]
  assign _GEN_100 = state ? _GEN_78 : _GEN_18; // @[Conditional.scala 39:67]
  assign _GEN_101 = state ? _GEN_79 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_102 = state ? _GEN_80 : _GEN_22; // @[Conditional.scala 39:67]
  assign _GEN_103 = state ? _GEN_81 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_104 = state ? _GEN_82 : _GEN_26; // @[Conditional.scala 39:67]
  assign _GEN_105 = state ? _GEN_83 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_106 = state ? _GEN_84 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_107 = state ? _GEN_85 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_108 = state ? _GEN_86 : _GEN_34; // @[Conditional.scala 39:67]
  assign _GEN_110 = state ? _GEN_88 : state; // @[Conditional.scala 39:67]
  assign _GEN_111 = _T_526 ? _GEN_47 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_112 = _T_526 ? _GEN_48 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_113 = _T_526 ? _GEN_49 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_114 = _T_526 ? _GEN_50 : _GEN_7; // @[Conditional.scala 40:58]
  assign _GEN_115 = _T_526 ? _GEN_51 : _GEN_9; // @[Conditional.scala 40:58]
  assign _GEN_116 = _T_526 ? _GEN_52 : _GEN_11; // @[Conditional.scala 40:58]
  assign _GEN_117 = _T_526 ? _GEN_53 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_118 = _T_526 ? _GEN_54 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_119 = _T_526 ? _GEN_55 : _GEN_17; // @[Conditional.scala 40:58]
  assign _GEN_120 = _T_526 ? _GEN_56 : _GEN_19; // @[Conditional.scala 40:58]
  assign _GEN_121 = _T_526 ? _GEN_57 : _GEN_21; // @[Conditional.scala 40:58]
  assign _GEN_122 = _T_526 ? _GEN_58 : _GEN_23; // @[Conditional.scala 40:58]
  assign _GEN_123 = _T_526 ? _GEN_59 : _GEN_25; // @[Conditional.scala 40:58]
  assign _GEN_124 = _T_526 ? _GEN_60 : _GEN_27; // @[Conditional.scala 40:58]
  assign _GEN_125 = _T_526 ? _GEN_61 : _GEN_29; // @[Conditional.scala 40:58]
  assign _GEN_126 = _T_526 ? _GEN_62 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_127 = _T_526 ? _GEN_63 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_128 = _T_526 ? _GEN_64 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_129 = _T_526 ? _GEN_65 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_130 = _T_526 ? _GEN_66 : _GEN_110; // @[Conditional.scala 40:58]
  assign _GEN_131 = _T_526 ? _GEN_42 : _GEN_89; // @[Conditional.scala 40:58]
  assign _GEN_132 = _T_526 ? _GEN_46 : _GEN_90; // @[Conditional.scala 40:58]
  assign _GEN_133 = _T_526 ? _GEN_0 : _GEN_91; // @[Conditional.scala 40:58]
  assign _GEN_134 = _T_526 ? _GEN_2 : _GEN_92; // @[Conditional.scala 40:58]
  assign _GEN_135 = _T_526 ? _GEN_4 : _GEN_93; // @[Conditional.scala 40:58]
  assign _GEN_136 = _T_526 ? _GEN_6 : _GEN_94; // @[Conditional.scala 40:58]
  assign _GEN_137 = _T_526 ? _GEN_8 : _GEN_95; // @[Conditional.scala 40:58]
  assign _GEN_138 = _T_526 ? _GEN_10 : _GEN_96; // @[Conditional.scala 40:58]
  assign _GEN_139 = _T_526 ? _GEN_12 : _GEN_97; // @[Conditional.scala 40:58]
  assign _GEN_140 = _T_526 ? _GEN_14 : _GEN_98; // @[Conditional.scala 40:58]
  assign _GEN_141 = _T_526 ? _GEN_16 : _GEN_99; // @[Conditional.scala 40:58]
  assign _GEN_142 = _T_526 ? _GEN_18 : _GEN_100; // @[Conditional.scala 40:58]
  assign _GEN_143 = _T_526 ? _GEN_20 : _GEN_101; // @[Conditional.scala 40:58]
  assign _GEN_144 = _T_526 ? _GEN_22 : _GEN_102; // @[Conditional.scala 40:58]
  assign _GEN_145 = _T_526 ? _GEN_24 : _GEN_103; // @[Conditional.scala 40:58]
  assign _GEN_146 = _T_526 ? _GEN_26 : _GEN_104; // @[Conditional.scala 40:58]
  assign _GEN_147 = _T_526 ? _GEN_28 : _GEN_105; // @[Conditional.scala 40:58]
  assign _GEN_148 = _T_526 ? _GEN_30 : _GEN_106; // @[Conditional.scala 40:58]
  assign _GEN_149 = _T_526 ? _GEN_32 : _GEN_107; // @[Conditional.scala 40:58]
  assign _GEN_150 = _T_526 ? _GEN_34 : _GEN_108; // @[Conditional.scala 40:58]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 733:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 111:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 722:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 722:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 722:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 722:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 722:21]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 722:21]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 722:21]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 722:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 722:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_8_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 722:21]
  assign io_Out_9_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_10_valid = out_valid_R_10; // @[HandShaking.scala 722:21]
  assign io_Out_10_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_11_valid = out_valid_R_11; // @[HandShaking.scala 722:21]
  assign io_Out_11_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_12_valid = out_valid_R_12; // @[HandShaking.scala 722:21]
  assign io_Out_12_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_12_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_13_valid = out_valid_R_13; // @[HandShaking.scala 722:21]
  assign io_Out_13_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_13_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_14_valid = out_valid_R_14; // @[HandShaking.scala 722:21]
  assign io_Out_14_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_14_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_15_valid = out_valid_R_15; // @[HandShaking.scala 722:21]
  assign io_Out_15_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_15_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_16_valid = out_valid_R_16; // @[HandShaking.scala 722:21]
  assign io_Out_16_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_16_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_Out_17_valid = out_valid_R_17; // @[HandShaking.scala 722:21]
  assign io_Out_17_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 106:27]
  assign io_Out_17_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 105:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 95:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 95:29]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_ready_R_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_ready_R_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_ready_R_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_ready_R_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_ready_R_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_ready_R_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_valid_R_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_valid_R_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_valid_R_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_valid_R_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_valid_R_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_valid_R_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_valid_R_16 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_valid_R_17 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_37[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_39[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  state = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_425) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_425) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_425) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_427) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_427) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_427) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_429) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_429) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_429) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_431) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_431) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_431) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_433) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_433) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_433) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_435) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_435) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_435) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_437) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_437) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_437) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_439) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_439) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_439) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_441) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_441) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_441) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_443) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_443) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_443) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_10 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_445) begin
          out_ready_R_10 <= io_Out_10_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_10 <= 1'h0;
          end else begin
            if (_T_445) begin
              out_ready_R_10 <= io_Out_10_ready;
            end
          end
        end else begin
          if (_T_445) begin
            out_ready_R_10 <= io_Out_10_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_11 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_447) begin
          out_ready_R_11 <= io_Out_11_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_11 <= 1'h0;
          end else begin
            if (_T_447) begin
              out_ready_R_11 <= io_Out_11_ready;
            end
          end
        end else begin
          if (_T_447) begin
            out_ready_R_11 <= io_Out_11_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_12 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_449) begin
          out_ready_R_12 <= io_Out_12_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_12 <= 1'h0;
          end else begin
            if (_T_449) begin
              out_ready_R_12 <= io_Out_12_ready;
            end
          end
        end else begin
          if (_T_449) begin
            out_ready_R_12 <= io_Out_12_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_13 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_451) begin
          out_ready_R_13 <= io_Out_13_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_13 <= 1'h0;
          end else begin
            if (_T_451) begin
              out_ready_R_13 <= io_Out_13_ready;
            end
          end
        end else begin
          if (_T_451) begin
            out_ready_R_13 <= io_Out_13_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_14 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_453) begin
          out_ready_R_14 <= io_Out_14_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_14 <= 1'h0;
          end else begin
            if (_T_453) begin
              out_ready_R_14 <= io_Out_14_ready;
            end
          end
        end else begin
          if (_T_453) begin
            out_ready_R_14 <= io_Out_14_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_15 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_455) begin
          out_ready_R_15 <= io_Out_15_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_15 <= 1'h0;
          end else begin
            if (_T_455) begin
              out_ready_R_15 <= io_Out_15_ready;
            end
          end
        end else begin
          if (_T_455) begin
            out_ready_R_15 <= io_Out_15_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_16 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_457) begin
          out_ready_R_16 <= io_Out_16_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_16 <= 1'h0;
          end else begin
            if (_T_457) begin
              out_ready_R_16 <= io_Out_16_ready;
            end
          end
        end else begin
          if (_T_457) begin
            out_ready_R_16 <= io_Out_16_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_17 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_459) begin
          out_ready_R_17 <= io_Out_17_ready;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            out_ready_R_17 <= 1'h0;
          end else begin
            if (_T_459) begin
              out_ready_R_17 <= io_Out_17_ready;
            end
          end
        end else begin
          if (_T_459) begin
            out_ready_R_17 <= io_Out_17_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_425) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_425) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_427) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_427) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_2 <= 1'h1;
        end else begin
          if (_T_429) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_429) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_3 <= 1'h1;
        end else begin
          if (_T_431) begin
            out_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_431) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_4 <= 1'h1;
        end else begin
          if (_T_433) begin
            out_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_433) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_5 <= 1'h1;
        end else begin
          if (_T_435) begin
            out_valid_R_5 <= 1'h0;
          end
        end
      end else begin
        if (_T_435) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_6 <= 1'h1;
        end else begin
          if (_T_437) begin
            out_valid_R_6 <= 1'h0;
          end
        end
      end else begin
        if (_T_437) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_7 <= 1'h1;
        end else begin
          if (_T_439) begin
            out_valid_R_7 <= 1'h0;
          end
        end
      end else begin
        if (_T_439) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_8 <= 1'h1;
        end else begin
          if (_T_441) begin
            out_valid_R_8 <= 1'h0;
          end
        end
      end else begin
        if (_T_441) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_9 <= 1'h1;
        end else begin
          if (_T_443) begin
            out_valid_R_9 <= 1'h0;
          end
        end
      end else begin
        if (_T_443) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_10 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_10 <= 1'h1;
        end else begin
          if (_T_445) begin
            out_valid_R_10 <= 1'h0;
          end
        end
      end else begin
        if (_T_445) begin
          out_valid_R_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_11 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_11 <= 1'h1;
        end else begin
          if (_T_447) begin
            out_valid_R_11 <= 1'h0;
          end
        end
      end else begin
        if (_T_447) begin
          out_valid_R_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_12 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_12 <= 1'h1;
        end else begin
          if (_T_449) begin
            out_valid_R_12 <= 1'h0;
          end
        end
      end else begin
        if (_T_449) begin
          out_valid_R_12 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_13 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_13 <= 1'h1;
        end else begin
          if (_T_451) begin
            out_valid_R_13 <= 1'h0;
          end
        end
      end else begin
        if (_T_451) begin
          out_valid_R_13 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_14 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_14 <= 1'h1;
        end else begin
          if (_T_453) begin
            out_valid_R_14 <= 1'h0;
          end
        end
      end else begin
        if (_T_453) begin
          out_valid_R_14 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_15 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_15 <= 1'h1;
        end else begin
          if (_T_455) begin
            out_valid_R_15 <= 1'h0;
          end
        end
      end else begin
        if (_T_455) begin
          out_valid_R_15 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_16 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_16 <= 1'h1;
        end else begin
          if (_T_457) begin
            out_valid_R_16 <= 1'h0;
          end
        end
      end else begin
        if (_T_457) begin
          out_valid_R_16 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_17 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          out_valid_R_17 <= 1'h1;
        end else begin
          if (_T_459) begin
            out_valid_R_17 <= 1'h0;
          end
        end
      end else begin
        if (_T_459) begin
          out_valid_R_17 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          mask_valid_R_0 <= 1'h1;
        end else begin
          if (_T_461) begin
            mask_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_461) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 10'h0;
    end else begin
      if (_T_515) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_515) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 10'h0;
    end else begin
      if (_T_516) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_516) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_515) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_516) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_515) begin
          predicate_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            if (_T_515) begin
              predicate_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_515) begin
            predicate_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_526) begin
        if (_T_516) begin
          predicate_valid_R_1 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            if (_T_516) begin
              predicate_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_516) begin
            predicate_valid_R_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_526) begin
        if (start) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_590) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module BasicBlockNoMaskFastNode_1(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [9:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [9:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [9:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [9:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [9:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
  reg [9:0] in_data_R_0_taskID; // @[BasicBlock.scala 988:46]
  reg [31:0] _RAND_0;
  reg  in_data_R_0_control; // @[BasicBlock.scala 988:46]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 989:52]
  reg [31:0] _RAND_2;
  reg [9:0] output_R_taskID; // @[BasicBlock.scala 991:25]
  reg [31:0] _RAND_3;
  reg  output_R_control; // @[BasicBlock.scala 991:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 992:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 992:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 992:49]
  reg [31:0] _RAND_7;
  reg  output_valid_R_3; // @[BasicBlock.scala 992:49]
  reg [31:0] _RAND_8;
  reg  output_valid_R_4; // @[BasicBlock.scala 992:49]
  reg [31:0] _RAND_9;
  reg  output_fire_R_0; // @[BasicBlock.scala 993:48]
  reg [31:0] _RAND_10;
  reg  output_fire_R_1; // @[BasicBlock.scala 993:48]
  reg [31:0] _RAND_11;
  reg  output_fire_R_2; // @[BasicBlock.scala 993:48]
  reg [31:0] _RAND_12;
  reg  output_fire_R_3; // @[BasicBlock.scala 993:48]
  reg [31:0] _RAND_13;
  reg  output_fire_R_4; // @[BasicBlock.scala 993:48]
  reg [31:0] _RAND_14;
  wire  _T_105; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_1; // @[BasicBlock.scala 998:36]
  wire  _GEN_2; // @[BasicBlock.scala 998:36]
  wire  _GEN_3; // @[BasicBlock.scala 998:36]
  wire [9:0] in_task_ID; // @[BasicBlock.scala 1005:34]
  wire  _T_107; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[BasicBlock.scala 1010:28]
  wire  _GEN_5; // @[BasicBlock.scala 1010:28]
  wire  _T_110; // @[Decoupled.scala 37:37]
  wire  _GEN_6; // @[BasicBlock.scala 1010:28]
  wire  _GEN_7; // @[BasicBlock.scala 1010:28]
  wire  _T_113; // @[Decoupled.scala 37:37]
  wire  _GEN_8; // @[BasicBlock.scala 1010:28]
  wire  _GEN_9; // @[BasicBlock.scala 1010:28]
  wire  _T_116; // @[Decoupled.scala 37:37]
  wire  _GEN_10; // @[BasicBlock.scala 1010:28]
  wire  _GEN_11; // @[BasicBlock.scala 1010:28]
  wire  _T_119; // @[Decoupled.scala 37:37]
  wire  _GEN_12; // @[BasicBlock.scala 1010:28]
  wire  _GEN_13; // @[BasicBlock.scala 1010:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 1027:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 1027:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 1027:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 1027:85]
  wire  out_fire_mask_4; // @[BasicBlock.scala 1027:85]
  reg  state; // @[BasicBlock.scala 1040:22]
  reg [31:0] _RAND_15;
  wire  _T_131; // @[Conditional.scala 37:30]
  wire  _GEN_14; // @[BasicBlock.scala 1045:43]
  wire  _GEN_15; // @[BasicBlock.scala 1045:43]
  wire  _GEN_16; // @[BasicBlock.scala 1045:43]
  wire  _GEN_17; // @[BasicBlock.scala 1045:43]
  wire  _GEN_18; // @[BasicBlock.scala 1045:43]
  wire  _GEN_19; // @[BasicBlock.scala 1045:43]
  wire  _T_138; // @[BasicBlock.scala 1066:35]
  wire  _T_139; // @[BasicBlock.scala 1066:35]
  wire  _T_140; // @[BasicBlock.scala 1066:35]
  wire  _T_141; // @[BasicBlock.scala 1066:35]
  wire  _GEN_20; // @[BasicBlock.scala 1066:41]
  wire [9:0] _GEN_21; // @[BasicBlock.scala 1066:41]
  wire  _GEN_22; // @[BasicBlock.scala 1066:41]
  wire  _GEN_23; // @[BasicBlock.scala 1066:41]
  wire  _GEN_24; // @[BasicBlock.scala 1066:41]
  wire  _GEN_25; // @[BasicBlock.scala 1066:41]
  wire  _GEN_26; // @[BasicBlock.scala 1066:41]
  wire  _GEN_27; // @[BasicBlock.scala 1066:41]
  wire  _GEN_28; // @[BasicBlock.scala 1066:41]
  wire  _GEN_29; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_32; // @[Conditional.scala 39:67]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 40:58]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire  _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire  _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  wire  _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  assign _T_105 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_105 ? io_predicateIn_0_bits_taskID : in_data_R_0_taskID; // @[BasicBlock.scala 998:36]
  assign _GEN_2 = _T_105 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 998:36]
  assign _GEN_3 = _T_105 ? 1'h1 : in_data_valid_R_0; // @[BasicBlock.scala 998:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 1005:34]
  assign _T_107 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_107 ? 1'h1 : output_fire_R_0; // @[BasicBlock.scala 1010:28]
  assign _GEN_5 = _T_107 ? 1'h0 : output_valid_R_0; // @[BasicBlock.scala 1010:28]
  assign _T_110 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_110 ? 1'h1 : output_fire_R_1; // @[BasicBlock.scala 1010:28]
  assign _GEN_7 = _T_110 ? 1'h0 : output_valid_R_1; // @[BasicBlock.scala 1010:28]
  assign _T_113 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_113 ? 1'h1 : output_fire_R_2; // @[BasicBlock.scala 1010:28]
  assign _GEN_9 = _T_113 ? 1'h0 : output_valid_R_2; // @[BasicBlock.scala 1010:28]
  assign _T_116 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 37:37]
  assign _GEN_10 = _T_116 ? 1'h1 : output_fire_R_3; // @[BasicBlock.scala 1010:28]
  assign _GEN_11 = _T_116 ? 1'h0 : output_valid_R_3; // @[BasicBlock.scala 1010:28]
  assign _T_119 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_119 ? 1'h1 : output_fire_R_4; // @[BasicBlock.scala 1010:28]
  assign _GEN_13 = _T_119 ? 1'h0 : output_valid_R_4; // @[BasicBlock.scala 1010:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_107; // @[BasicBlock.scala 1027:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_110; // @[BasicBlock.scala 1027:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_113; // @[BasicBlock.scala 1027:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_116; // @[BasicBlock.scala 1027:85]
  assign out_fire_mask_4 = output_fire_R_4 | _T_119; // @[BasicBlock.scala 1027:85]
  assign _T_131 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_14 = in_data_valid_R_0 ? 1'h1 : _GEN_5; // @[BasicBlock.scala 1045:43]
  assign _GEN_15 = in_data_valid_R_0 ? 1'h1 : _GEN_7; // @[BasicBlock.scala 1045:43]
  assign _GEN_16 = in_data_valid_R_0 ? 1'h1 : _GEN_9; // @[BasicBlock.scala 1045:43]
  assign _GEN_17 = in_data_valid_R_0 ? 1'h1 : _GEN_11; // @[BasicBlock.scala 1045:43]
  assign _GEN_18 = in_data_valid_R_0 ? 1'h1 : _GEN_13; // @[BasicBlock.scala 1045:43]
  assign _GEN_19 = in_data_valid_R_0 ? 1'h1 : state; // @[BasicBlock.scala 1045:43]
  assign _T_138 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 1066:35]
  assign _T_139 = _T_138 & out_fire_mask_2; // @[BasicBlock.scala 1066:35]
  assign _T_140 = _T_139 & out_fire_mask_3; // @[BasicBlock.scala 1066:35]
  assign _T_141 = _T_140 & out_fire_mask_4; // @[BasicBlock.scala 1066:35]
  assign _GEN_20 = _T_141 ? 1'h0 : _GEN_2; // @[BasicBlock.scala 1066:41]
  assign _GEN_21 = _T_141 ? 10'h0 : _GEN_1; // @[BasicBlock.scala 1066:41]
  assign _GEN_22 = _T_141 ? 1'h0 : _GEN_3; // @[BasicBlock.scala 1066:41]
  assign _GEN_23 = _T_141 ? 1'h0 : _GEN_4; // @[BasicBlock.scala 1066:41]
  assign _GEN_24 = _T_141 ? 1'h0 : _GEN_6; // @[BasicBlock.scala 1066:41]
  assign _GEN_25 = _T_141 ? 1'h0 : _GEN_8; // @[BasicBlock.scala 1066:41]
  assign _GEN_26 = _T_141 ? 1'h0 : _GEN_10; // @[BasicBlock.scala 1066:41]
  assign _GEN_27 = _T_141 ? 1'h0 : _GEN_12; // @[BasicBlock.scala 1066:41]
  assign _GEN_28 = _T_141 ? 1'h0 : state; // @[BasicBlock.scala 1066:41]
  assign _GEN_29 = state ? _GEN_20 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_30 = state ? _GEN_21 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_31 = state ? _GEN_22 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_32 = state ? _GEN_23 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_33 = state ? _GEN_24 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_25 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_26 : _GEN_10; // @[Conditional.scala 39:67]
  assign _GEN_36 = state ? _GEN_27 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_28 : state; // @[Conditional.scala 39:67]
  assign _GEN_38 = _T_131 ? _GEN_14 : _GEN_5; // @[Conditional.scala 40:58]
  assign _GEN_39 = _T_131 ? _GEN_15 : _GEN_7; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_131 ? _GEN_16 : _GEN_9; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_131 ? _GEN_17 : _GEN_11; // @[Conditional.scala 40:58]
  assign _GEN_42 = _T_131 ? _GEN_18 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_131 ? _GEN_19 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_131 ? _GEN_2 : _GEN_29; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_131 ? _GEN_1 : _GEN_30; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_131 ? _GEN_3 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_131 ? _GEN_4 : _GEN_32; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_131 ? _GEN_6 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_131 ? _GEN_8 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_131 ? _GEN_10 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_131 ? _GEN_12 : _GEN_36; // @[Conditional.scala 40:58]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 997:29]
  assign io_Out_0_valid = output_valid_R_0; // @[BasicBlock.scala 1019:21]
  assign io_Out_0_bits_taskID = output_R_taskID; // @[BasicBlock.scala 1018:20]
  assign io_Out_1_valid = output_valid_R_1; // @[BasicBlock.scala 1019:21]
  assign io_Out_1_bits_taskID = output_R_taskID; // @[BasicBlock.scala 1018:20]
  assign io_Out_2_valid = output_valid_R_2; // @[BasicBlock.scala 1019:21]
  assign io_Out_2_bits_taskID = output_R_taskID; // @[BasicBlock.scala 1018:20]
  assign io_Out_2_bits_control = output_R_control; // @[BasicBlock.scala 1018:20]
  assign io_Out_3_valid = output_valid_R_3; // @[BasicBlock.scala 1019:21]
  assign io_Out_3_bits_taskID = output_R_taskID; // @[BasicBlock.scala 1018:20]
  assign io_Out_3_bits_control = output_R_control; // @[BasicBlock.scala 1018:20]
  assign io_Out_4_valid = output_valid_R_4; // @[BasicBlock.scala 1019:21]
  assign io_Out_4_bits_taskID = output_R_taskID; // @[BasicBlock.scala 1018:20]
  assign io_Out_4_bits_control = output_R_control; // @[BasicBlock.scala 1018:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  output_R_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      in_data_R_0_taskID <= 10'h0;
    end else begin
      if (_T_131) begin
        if (_T_105) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            in_data_R_0_taskID <= 10'h0;
          end else begin
            if (_T_105) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_105) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_105) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_105) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_105) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_105) begin
          in_data_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            if (_T_105) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_105) begin
            in_data_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 10'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_R_control <= 1'h0;
    end else begin
      output_R_control <= in_data_R_0_control;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (in_data_valid_R_0) begin
          output_valid_R_0 <= 1'h1;
        end else begin
          if (_T_107) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_107) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (in_data_valid_R_0) begin
          output_valid_R_1 <= 1'h1;
        end else begin
          if (_T_110) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_110) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (in_data_valid_R_0) begin
          output_valid_R_2 <= 1'h1;
        end else begin
          if (_T_113) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_113) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (in_data_valid_R_0) begin
          output_valid_R_3 <= 1'h1;
        end else begin
          if (_T_116) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_116) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (in_data_valid_R_0) begin
          output_valid_R_4 <= 1'h1;
        end else begin
          if (_T_119) begin
            output_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_119) begin
          output_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_107) begin
          output_fire_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            if (_T_107) begin
              output_fire_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_107) begin
            output_fire_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_110) begin
          output_fire_R_1 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            if (_T_110) begin
              output_fire_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_110) begin
            output_fire_R_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_113) begin
          output_fire_R_2 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            if (_T_113) begin
              output_fire_R_2 <= 1'h1;
            end
          end
        end else begin
          if (_T_113) begin
            output_fire_R_2 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_116) begin
          output_fire_R_3 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            if (_T_116) begin
              output_fire_R_3 <= 1'h1;
            end
          end
        end else begin
          if (_T_116) begin
            output_fire_R_3 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else begin
      if (_T_131) begin
        if (_T_119) begin
          output_fire_R_4 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            output_fire_R_4 <= 1'h0;
          end else begin
            if (_T_119) begin
              output_fire_R_4 <= 1'h1;
            end
          end
        end else begin
          if (_T_119) begin
            output_fire_R_4 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_131) begin
        if (in_data_valid_R_0) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_141) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UBranchNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_142; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_145; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_5;
  wire  _T_156; // @[Conditional.scala 37:30]
  wire  _GEN_6; // @[BranchNode.scala 611:46]
  wire  _GEN_7; // @[BranchNode.scala 611:46]
  wire  _T_168; // @[HandShaking.scala 656:24]
  wire  _T_170; // @[HandShaking.scala 656:24]
  wire  _T_171; // @[HandShaking.scala 656:50]
  wire  _T_173; // @[HandShaking.scala 656:50]
  wire  _T_174; // @[HandShaking.scala 656:29]
  wire  _GEN_8; // @[BranchNode.scala 631:26]
  wire  _GEN_9; // @[BranchNode.scala 631:26]
  wire  _GEN_10; // @[BranchNode.scala 631:26]
  wire  _GEN_11; // @[BranchNode.scala 631:26]
  wire [9:0] _GEN_12; // @[BranchNode.scala 631:26]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_21; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_23; // @[Conditional.scala 40:58]
  assign _T_142 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_142 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_142 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_145 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_145 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_145 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_145 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_156 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_6 = enable_valid_R ? 1'h1 : state; // @[BranchNode.scala 611:46]
  assign _GEN_7 = enable_valid_R ? 1'h1 : _GEN_1; // @[BranchNode.scala 611:46]
  assign _T_168 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_170 = _T_168 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_171 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_173 = _T_171 == 1'h0; // @[HandShaking.scala 656:50]
  assign _T_174 = _T_170 | _T_173; // @[HandShaking.scala 656:29]
  assign _GEN_8 = _T_174 ? 1'h0 : state; // @[BranchNode.scala 631:26]
  assign _GEN_9 = _T_174 ? 1'h0 : _GEN_0; // @[BranchNode.scala 631:26]
  assign _GEN_10 = _T_174 ? 1'h0 : _GEN_2; // @[BranchNode.scala 631:26]
  assign _GEN_11 = _T_174 ? 1'h0 : _GEN_3; // @[BranchNode.scala 631:26]
  assign _GEN_12 = _T_174 ? 10'h0 : _GEN_4; // @[BranchNode.scala 631:26]
  assign _GEN_13 = state ? _GEN_8 : state; // @[Conditional.scala 39:67]
  assign _GEN_14 = state ? _GEN_9 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_11 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_12 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_156 ? _GEN_6 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_156 ? _GEN_7 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_156 ? _GEN_0 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_156 ? _GEN_2 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_156 ? _GEN_3 : _GEN_16; // @[Conditional.scala 40:58]
  assign _GEN_23 = _T_156 ? _GEN_4 : _GEN_17; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 606:20]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 606:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_145) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_145) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_142) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_142) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_142) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_142) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_142) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module PhiFastNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [9:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [9:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data
);
  reg [9:0] in_data_R_0_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_0;
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [9:0] in_data_R_1_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_5;
  reg [9:0] enable_R_taskID; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_6;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_7;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_8;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_9;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_10;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_12;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_13;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  wire  _T_172; // @[Decoupled.scala 37:37]
  wire [1:0] _GEN_1; // @[PhiNode.scala 215:24]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_175; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[PhiNode.scala 222:26]
  wire  _GEN_4; // @[PhiNode.scala 222:26]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_178; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[PhiNode.scala 230:29]
  wire [31:0] _GEN_8; // @[PhiNode.scala 230:29]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_181; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[PhiNode.scala 230:29]
  wire [31:0] _GEN_12; // @[PhiNode.scala 230:29]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [9:0] task_input; // @[PhiNode.scala 250:43]
  wire [9:0] _GEN_18; // @[PhiNode.scala 253:20]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_195; // @[Decoupled.scala 37:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_198; // @[Decoupled.scala 37:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_15;
  wire  _T_204; // @[Conditional.scala 37:30]
  wire  _T_205; // @[PhiNode.scala 268:37]
  wire  _T_206; // @[PhiNode.scala 277:27]
  wire [1:0] _GEN_24; // @[PhiNode.scala 279:32]
  wire  _GEN_25; // @[PhiNode.scala 277:46]
  wire  _GEN_26; // @[PhiNode.scala 277:46]
  wire [1:0] _GEN_27; // @[PhiNode.scala 277:46]
  wire  _T_209; // @[Conditional.scala 37:30]
  wire  _T_210; // @[PhiNode.scala 299:31]
  wire [31:0] _GEN_28; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_29; // @[PhiNode.scala 299:37]
  wire [31:0] _GEN_31; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_32; // @[PhiNode.scala 299:37]
  wire  _GEN_34; // @[PhiNode.scala 299:37]
  wire  _GEN_35; // @[PhiNode.scala 299:37]
  wire [1:0] _GEN_36; // @[PhiNode.scala 299:37]
  wire  _GEN_37; // @[PhiNode.scala 299:37]
  wire  _GEN_38; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_39; // @[PhiNode.scala 299:37]
  wire  _GEN_40; // @[PhiNode.scala 299:37]
  wire  _GEN_41; // @[PhiNode.scala 299:37]
  wire  _GEN_42; // @[PhiNode.scala 299:37]
  wire [1:0] _GEN_43; // @[PhiNode.scala 299:37]
  wire  _T_232; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_60; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_64; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_66; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_67; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_69; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_72; // @[Conditional.scala 39:67]
  wire  _GEN_73; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_74; // @[Conditional.scala 39:67]
  wire  _GEN_75; // @[Conditional.scala 39:67]
  wire  _GEN_76; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_77; // @[Conditional.scala 39:67]
  wire  _GEN_78; // @[Conditional.scala 39:67]
  wire  _GEN_79; // @[Conditional.scala 39:67]
  wire  _GEN_80; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_81; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_82; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_83; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_85; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_86; // @[Conditional.scala 39:67]
  wire  _GEN_88; // @[Conditional.scala 39:67]
  wire  _GEN_89; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_90; // @[Conditional.scala 39:67]
  wire  _GEN_91; // @[Conditional.scala 39:67]
  wire  _GEN_92; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_93; // @[Conditional.scala 39:67]
  wire  _GEN_94; // @[Conditional.scala 39:67]
  wire  _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_96; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_97; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_98; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_102; // @[Conditional.scala 39:67]
  wire  _GEN_104; // @[Conditional.scala 40:58]
  wire  _GEN_105; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_106; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_107; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_108; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_110; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_111; // @[Conditional.scala 40:58]
  wire  _GEN_113; // @[Conditional.scala 40:58]
  wire  _GEN_114; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_115; // @[Conditional.scala 40:58]
  wire  _GEN_116; // @[Conditional.scala 40:58]
  wire  _GEN_117; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_118; // @[Conditional.scala 40:58]
  wire  _GEN_119; // @[Conditional.scala 40:58]
  wire  _GEN_120; // @[Conditional.scala 40:58]
  wire  _GEN_121; // @[Conditional.scala 40:58]
  assign _T_172 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_172 ? io_Mask_bits : mask_R; // @[PhiNode.scala 215:24]
  assign _GEN_2 = _T_172 ? 1'h1 : mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_175 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_175 ? io_enable_bits_taskID : enable_R_taskID; // @[PhiNode.scala 222:26]
  assign _GEN_4 = _T_175 ? io_enable_bits_control : enable_R_control; // @[PhiNode.scala 222:26]
  assign _GEN_5 = _T_175 ? 1'h1 : enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_178 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_178 ? io_InData_0_bits_taskID : in_data_R_0_taskID; // @[PhiNode.scala 230:29]
  assign _GEN_8 = _T_178 ? 32'h0 : in_data_R_0_data; // @[PhiNode.scala 230:29]
  assign _GEN_9 = _T_178 ? 1'h1 : in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_181 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_181 ? io_InData_1_bits_taskID : in_data_R_1_taskID; // @[PhiNode.scala 230:29]
  assign _GEN_12 = _T_181 ? io_InData_1_bits_data : in_data_R_1_data; // @[PhiNode.scala 230:29]
  assign _GEN_13 = _T_181 ? 1'h1 : in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign sel = mask_R[1]; // @[CircuitMath.scala 30:8]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[PhiNode.scala 250:43]
  assign _GEN_18 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 253:20]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_195 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_20 = _T_195 ? 1'h1 : fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_195 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_198 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_22 = _T_198 ? 1'h1 : fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_198 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_195; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_198; // @[PhiNode.scala 265:74]
  assign _T_204 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_205 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_206 = enable_valid_R & _T_205; // @[PhiNode.scala 277:27]
  assign _GEN_24 = enable_R_control ? 2'h1 : 2'h2; // @[PhiNode.scala 279:32]
  assign _GEN_25 = _T_206 ? 1'h1 : _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_26 = _T_206 ? 1'h1 : _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_27 = _T_206 ? _GEN_24 : state; // @[PhiNode.scala 277:46]
  assign _T_209 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_210 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _GEN_28 = _T_210 ? 32'h0 : _GEN_8; // @[PhiNode.scala 299:37]
  assign _GEN_29 = _T_210 ? 10'h0 : _GEN_7; // @[PhiNode.scala 299:37]
  assign _GEN_31 = _T_210 ? 32'h0 : _GEN_12; // @[PhiNode.scala 299:37]
  assign _GEN_32 = _T_210 ? 10'h0 : _GEN_11; // @[PhiNode.scala 299:37]
  assign _GEN_34 = _T_210 ? 1'h0 : _GEN_9; // @[PhiNode.scala 299:37]
  assign _GEN_35 = _T_210 ? 1'h0 : _GEN_13; // @[PhiNode.scala 299:37]
  assign _GEN_36 = _T_210 ? 2'h0 : _GEN_1; // @[PhiNode.scala 299:37]
  assign _GEN_37 = _T_210 ? 1'h0 : _GEN_2; // @[PhiNode.scala 299:37]
  assign _GEN_38 = _T_210 ? 1'h0 : _GEN_4; // @[PhiNode.scala 299:37]
  assign _GEN_39 = _T_210 ? 10'h0 : _GEN_3; // @[PhiNode.scala 299:37]
  assign _GEN_40 = _T_210 ? 1'h0 : _GEN_5; // @[PhiNode.scala 299:37]
  assign _GEN_41 = _T_210 ? 1'h0 : _GEN_20; // @[PhiNode.scala 299:37]
  assign _GEN_42 = _T_210 ? 1'h0 : _GEN_22; // @[PhiNode.scala 299:37]
  assign _GEN_43 = _T_210 ? 2'h0 : state; // @[PhiNode.scala 299:37]
  assign _T_232 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_60 = _T_232 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_64 = _T_232 ? task_input : _GEN_18; // @[Conditional.scala 39:67]
  assign _GEN_66 = _T_232 ? _GEN_28 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_67 = _T_232 ? _GEN_29 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_69 = _T_232 ? _GEN_31 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_70 = _T_232 ? _GEN_32 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_72 = _T_232 ? _GEN_34 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_73 = _T_232 ? _GEN_35 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_74 = _T_232 ? _GEN_36 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_75 = _T_232 ? _GEN_37 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_76 = _T_232 ? _GEN_38 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_77 = _T_232 ? _GEN_39 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_78 = _T_232 ? _GEN_40 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_79 = _T_232 ? _GEN_41 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_80 = _T_232 ? _GEN_42 : _GEN_22; // @[Conditional.scala 39:67]
  assign _GEN_81 = _T_232 ? _GEN_43 : state; // @[Conditional.scala 39:67]
  assign _GEN_82 = _T_209 ? _GEN_28 : _GEN_66; // @[Conditional.scala 39:67]
  assign _GEN_83 = _T_209 ? _GEN_29 : _GEN_67; // @[Conditional.scala 39:67]
  assign _GEN_85 = _T_209 ? _GEN_31 : _GEN_69; // @[Conditional.scala 39:67]
  assign _GEN_86 = _T_209 ? _GEN_32 : _GEN_70; // @[Conditional.scala 39:67]
  assign _GEN_88 = _T_209 ? _GEN_34 : _GEN_72; // @[Conditional.scala 39:67]
  assign _GEN_89 = _T_209 ? _GEN_35 : _GEN_73; // @[Conditional.scala 39:67]
  assign _GEN_90 = _T_209 ? _GEN_36 : _GEN_74; // @[Conditional.scala 39:67]
  assign _GEN_91 = _T_209 ? _GEN_37 : _GEN_75; // @[Conditional.scala 39:67]
  assign _GEN_92 = _T_209 ? _GEN_38 : _GEN_76; // @[Conditional.scala 39:67]
  assign _GEN_93 = _T_209 ? _GEN_39 : _GEN_77; // @[Conditional.scala 39:67]
  assign _GEN_94 = _T_209 ? _GEN_40 : _GEN_78; // @[Conditional.scala 39:67]
  assign _GEN_95 = _T_209 ? _GEN_41 : _GEN_79; // @[Conditional.scala 39:67]
  assign _GEN_96 = _T_209 ? _GEN_42 : _GEN_80; // @[Conditional.scala 39:67]
  assign _GEN_97 = _T_209 ? _GEN_43 : _GEN_81; // @[Conditional.scala 39:67]
  assign _GEN_98 = _T_209 ? _GEN_19 : _GEN_60; // @[Conditional.scala 39:67]
  assign _GEN_102 = _T_209 ? _GEN_18 : _GEN_64; // @[Conditional.scala 39:67]
  assign _GEN_104 = _T_204 ? _GEN_25 : _GEN_21; // @[Conditional.scala 40:58]
  assign _GEN_105 = _T_204 ? _GEN_26 : _GEN_23; // @[Conditional.scala 40:58]
  assign _GEN_106 = _T_204 ? _GEN_27 : _GEN_97; // @[Conditional.scala 40:58]
  assign _GEN_107 = _T_204 ? _GEN_8 : _GEN_82; // @[Conditional.scala 40:58]
  assign _GEN_108 = _T_204 ? _GEN_7 : _GEN_83; // @[Conditional.scala 40:58]
  assign _GEN_110 = _T_204 ? _GEN_12 : _GEN_85; // @[Conditional.scala 40:58]
  assign _GEN_111 = _T_204 ? _GEN_11 : _GEN_86; // @[Conditional.scala 40:58]
  assign _GEN_113 = _T_204 ? _GEN_9 : _GEN_88; // @[Conditional.scala 40:58]
  assign _GEN_114 = _T_204 ? _GEN_13 : _GEN_89; // @[Conditional.scala 40:58]
  assign _GEN_115 = _T_204 ? _GEN_1 : _GEN_90; // @[Conditional.scala 40:58]
  assign _GEN_116 = _T_204 ? _GEN_2 : _GEN_91; // @[Conditional.scala 40:58]
  assign _GEN_117 = _T_204 ? _GEN_4 : _GEN_92; // @[Conditional.scala 40:58]
  assign _GEN_118 = _T_204 ? _GEN_3 : _GEN_93; // @[Conditional.scala 40:58]
  assign _GEN_119 = _T_204 ? _GEN_5 : _GEN_94; // @[Conditional.scala 40:58]
  assign _GEN_120 = _T_204 ? _GEN_20 : _GEN_95; // @[Conditional.scala 40:58]
  assign _GEN_121 = _T_204 ? _GEN_22 : _GEN_96; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_204 ? _GEN_19 : _GEN_98; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_taskID = _T_204 ? _GEN_18 : _GEN_102; // @[PhiNode.scala 253:20 PhiNode.scala 326:44]
  assign io_Out_1_bits_data = _T_204 ? _GEN_19 : _GEN_98; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enable_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enable_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mask_R = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      in_data_R_0_taskID <= 10'h0;
    end else begin
      if (_T_204) begin
        if (_T_178) begin
          in_data_R_0_taskID <= io_InData_0_bits_taskID;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            in_data_R_0_taskID <= 10'h0;
          end else begin
            if (_T_178) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              in_data_R_0_taskID <= 10'h0;
            end else begin
              if (_T_178) begin
                in_data_R_0_taskID <= io_InData_0_bits_taskID;
              end
            end
          end else begin
            if (_T_178) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_204) begin
        if (_T_178) begin
          in_data_R_0_data <= 32'h0;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_178) begin
              in_data_R_0_data <= 32'h0;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_178) begin
                in_data_R_0_data <= 32'h0;
              end
            end
          end else begin
            if (_T_178) begin
              in_data_R_0_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 10'h0;
    end else begin
      if (_T_204) begin
        if (_T_181) begin
          in_data_R_1_taskID <= io_InData_1_bits_taskID;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            in_data_R_1_taskID <= 10'h0;
          end else begin
            if (_T_181) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              in_data_R_1_taskID <= 10'h0;
            end else begin
              if (_T_181) begin
                in_data_R_1_taskID <= io_InData_1_bits_taskID;
              end
            end
          end else begin
            if (_T_181) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_204) begin
        if (_T_181) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_181) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_181) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_181) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_178) begin
          in_data_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            if (_T_178) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              if (_T_178) begin
                in_data_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_178) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_181) begin
          in_data_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            if (_T_181) begin
              in_data_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              if (_T_181) begin
                in_data_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_181) begin
              in_data_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_204) begin
        if (_T_175) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_175) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_175) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_175) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_175) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_175) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_175) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_175) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_175) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_175) begin
              enable_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_175) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_175) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_204) begin
        if (_T_172) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_172) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_172) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_172) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_172) begin
          mask_valid_R <= 1'h1;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            mask_valid_R <= 1'h0;
          end else begin
            if (_T_172) begin
              mask_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              mask_valid_R <= 1'h0;
            end else begin
              if (_T_172) begin
                mask_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_172) begin
              mask_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_206) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_195) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_195) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_206) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_198) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_198) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_195) begin
          fire_R_0 <= 1'h1;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            fire_R_0 <= 1'h0;
          end else begin
            if (_T_195) begin
              fire_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              fire_R_0 <= 1'h0;
            end else begin
              if (_T_195) begin
                fire_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_195) begin
              fire_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_204) begin
        if (_T_198) begin
          fire_R_1 <= 1'h1;
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            fire_R_1 <= 1'h0;
          end else begin
            if (_T_198) begin
              fire_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              fire_R_1 <= 1'h0;
            end else begin
              if (_T_198) begin
                fire_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_198) begin
              fire_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_204) begin
        if (_T_206) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_209) begin
          if (_T_210) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_232) begin
            if (_T_210) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module UBranchNode_1(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_142; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_145; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_5;
  wire  _T_156; // @[Conditional.scala 37:30]
  wire  _GEN_6; // @[BranchNode.scala 611:46]
  wire  _GEN_7; // @[BranchNode.scala 611:46]
  wire  _T_168; // @[HandShaking.scala 656:24]
  wire  _T_170; // @[HandShaking.scala 656:24]
  wire  _T_171; // @[HandShaking.scala 656:50]
  wire  _T_173; // @[HandShaking.scala 656:50]
  wire  _T_174; // @[HandShaking.scala 656:29]
  wire  _GEN_8; // @[BranchNode.scala 631:26]
  wire  _GEN_9; // @[BranchNode.scala 631:26]
  wire  _GEN_10; // @[BranchNode.scala 631:26]
  wire  _GEN_11; // @[BranchNode.scala 631:26]
  wire [9:0] _GEN_12; // @[BranchNode.scala 631:26]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_21; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_23; // @[Conditional.scala 40:58]
  assign _T_142 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_142 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_142 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_145 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_145 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_145 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_145 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_156 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_6 = enable_valid_R ? 1'h1 : state; // @[BranchNode.scala 611:46]
  assign _GEN_7 = enable_valid_R ? 1'h1 : _GEN_1; // @[BranchNode.scala 611:46]
  assign _T_168 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_170 = _T_168 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_171 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_173 = _T_171 == 1'h0; // @[HandShaking.scala 656:50]
  assign _T_174 = _T_170 | _T_173; // @[HandShaking.scala 656:29]
  assign _GEN_8 = _T_174 ? 1'h0 : state; // @[BranchNode.scala 631:26]
  assign _GEN_9 = _T_174 ? 1'h0 : _GEN_0; // @[BranchNode.scala 631:26]
  assign _GEN_10 = _T_174 ? 1'h0 : _GEN_2; // @[BranchNode.scala 631:26]
  assign _GEN_11 = _T_174 ? 1'h0 : _GEN_3; // @[BranchNode.scala 631:26]
  assign _GEN_12 = _T_174 ? 10'h0 : _GEN_4; // @[BranchNode.scala 631:26]
  assign _GEN_13 = state ? _GEN_8 : state; // @[Conditional.scala 39:67]
  assign _GEN_14 = state ? _GEN_9 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_11 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_12 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_156 ? _GEN_6 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_156 ? _GEN_7 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_156 ? _GEN_0 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_156 ? _GEN_2 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_156 ? _GEN_3 : _GEN_16; // @[Conditional.scala 40:58]
  assign _GEN_23 = _T_156 ? _GEN_4 : _GEN_17; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 606:20]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 606:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_145) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_145) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_142) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_142) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_142) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_142) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_142) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UBranchNode_2(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_142; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_145; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_5;
  wire  _T_156; // @[Conditional.scala 37:30]
  wire  _GEN_6; // @[BranchNode.scala 611:46]
  wire  _GEN_7; // @[BranchNode.scala 611:46]
  wire  _T_168; // @[HandShaking.scala 656:24]
  wire  _T_170; // @[HandShaking.scala 656:24]
  wire  _T_171; // @[HandShaking.scala 656:50]
  wire  _T_173; // @[HandShaking.scala 656:50]
  wire  _T_174; // @[HandShaking.scala 656:29]
  wire  _GEN_8; // @[BranchNode.scala 631:26]
  wire  _GEN_9; // @[BranchNode.scala 631:26]
  wire  _GEN_10; // @[BranchNode.scala 631:26]
  wire  _GEN_11; // @[BranchNode.scala 631:26]
  wire [9:0] _GEN_12; // @[BranchNode.scala 631:26]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_21; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_23; // @[Conditional.scala 40:58]
  assign _T_142 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_142 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_142 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_145 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_145 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_145 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_145 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_156 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_6 = enable_valid_R ? 1'h1 : state; // @[BranchNode.scala 611:46]
  assign _GEN_7 = enable_valid_R ? 1'h1 : _GEN_1; // @[BranchNode.scala 611:46]
  assign _T_168 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_170 = _T_168 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_171 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_173 = _T_171 == 1'h0; // @[HandShaking.scala 656:50]
  assign _T_174 = _T_170 | _T_173; // @[HandShaking.scala 656:29]
  assign _GEN_8 = _T_174 ? 1'h0 : state; // @[BranchNode.scala 631:26]
  assign _GEN_9 = _T_174 ? 1'h0 : _GEN_0; // @[BranchNode.scala 631:26]
  assign _GEN_10 = _T_174 ? 1'h0 : _GEN_2; // @[BranchNode.scala 631:26]
  assign _GEN_11 = _T_174 ? 1'h0 : _GEN_3; // @[BranchNode.scala 631:26]
  assign _GEN_12 = _T_174 ? 10'h0 : _GEN_4; // @[BranchNode.scala 631:26]
  assign _GEN_13 = state ? _GEN_8 : state; // @[Conditional.scala 39:67]
  assign _GEN_14 = state ? _GEN_9 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_11 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_12 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_156 ? _GEN_6 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_156 ? _GEN_7 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_156 ? _GEN_0 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_156 ? _GEN_2 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_156 ? _GEN_3 : _GEN_16; // @[Conditional.scala 40:58]
  assign _GEN_23 = _T_156 ? _GEN_4 : _GEN_17; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 606:20]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 606:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_145) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_145) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_142) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_142) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_142) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_142) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_142) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module PhiFastNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [9:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [9:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data
);
  reg [9:0] in_data_R_0_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_0;
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [9:0] in_data_R_1_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_5;
  reg [9:0] enable_R_taskID; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_6;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_7;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_8;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_9;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_10;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_12;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_13;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  wire  _T_172; // @[Decoupled.scala 37:37]
  wire [1:0] _GEN_1; // @[PhiNode.scala 215:24]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_175; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[PhiNode.scala 222:26]
  wire  _GEN_4; // @[PhiNode.scala 222:26]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_178; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[PhiNode.scala 230:29]
  wire [31:0] _GEN_8; // @[PhiNode.scala 230:29]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_181; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[PhiNode.scala 230:29]
  wire [31:0] _GEN_12; // @[PhiNode.scala 230:29]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_183; // @[Bitwise.scala 109:18]
  wire  _T_184; // @[Bitwise.scala 109:44]
  wire [1:0] _T_185; // @[Cat.scala 30:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [9:0] task_input; // @[PhiNode.scala 250:43]
  wire [9:0] _GEN_18; // @[PhiNode.scala 253:20]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_198; // @[Decoupled.scala 37:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_201; // @[Decoupled.scala 37:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_15;
  wire  _T_207; // @[Conditional.scala 37:30]
  wire  _T_208; // @[PhiNode.scala 268:37]
  wire  _T_209; // @[PhiNode.scala 277:27]
  wire [1:0] _GEN_24; // @[PhiNode.scala 279:32]
  wire  _GEN_25; // @[PhiNode.scala 277:46]
  wire  _GEN_26; // @[PhiNode.scala 277:46]
  wire [1:0] _GEN_27; // @[PhiNode.scala 277:46]
  wire  _T_212; // @[Conditional.scala 37:30]
  wire  _T_213; // @[PhiNode.scala 299:31]
  wire [31:0] _GEN_28; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_29; // @[PhiNode.scala 299:37]
  wire [31:0] _GEN_31; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_32; // @[PhiNode.scala 299:37]
  wire  _GEN_34; // @[PhiNode.scala 299:37]
  wire  _GEN_35; // @[PhiNode.scala 299:37]
  wire [1:0] _GEN_36; // @[PhiNode.scala 299:37]
  wire  _GEN_37; // @[PhiNode.scala 299:37]
  wire  _GEN_38; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_39; // @[PhiNode.scala 299:37]
  wire  _GEN_40; // @[PhiNode.scala 299:37]
  wire  _GEN_41; // @[PhiNode.scala 299:37]
  wire  _GEN_42; // @[PhiNode.scala 299:37]
  wire [1:0] _GEN_43; // @[PhiNode.scala 299:37]
  wire  _T_235; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_60; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_64; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_66; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_67; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_69; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_72; // @[Conditional.scala 39:67]
  wire  _GEN_73; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_74; // @[Conditional.scala 39:67]
  wire  _GEN_75; // @[Conditional.scala 39:67]
  wire  _GEN_76; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_77; // @[Conditional.scala 39:67]
  wire  _GEN_78; // @[Conditional.scala 39:67]
  wire  _GEN_79; // @[Conditional.scala 39:67]
  wire  _GEN_80; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_81; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_82; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_83; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_85; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_86; // @[Conditional.scala 39:67]
  wire  _GEN_88; // @[Conditional.scala 39:67]
  wire  _GEN_89; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_90; // @[Conditional.scala 39:67]
  wire  _GEN_91; // @[Conditional.scala 39:67]
  wire  _GEN_92; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_93; // @[Conditional.scala 39:67]
  wire  _GEN_94; // @[Conditional.scala 39:67]
  wire  _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_96; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_97; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_98; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_102; // @[Conditional.scala 39:67]
  wire  _GEN_104; // @[Conditional.scala 40:58]
  wire  _GEN_105; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_106; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_107; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_108; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_110; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_111; // @[Conditional.scala 40:58]
  wire  _GEN_113; // @[Conditional.scala 40:58]
  wire  _GEN_114; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_115; // @[Conditional.scala 40:58]
  wire  _GEN_116; // @[Conditional.scala 40:58]
  wire  _GEN_117; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_118; // @[Conditional.scala 40:58]
  wire  _GEN_119; // @[Conditional.scala 40:58]
  wire  _GEN_120; // @[Conditional.scala 40:58]
  wire  _GEN_121; // @[Conditional.scala 40:58]
  assign _T_172 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_172 ? io_Mask_bits : mask_R; // @[PhiNode.scala 215:24]
  assign _GEN_2 = _T_172 ? 1'h1 : mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_175 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_175 ? io_enable_bits_taskID : enable_R_taskID; // @[PhiNode.scala 222:26]
  assign _GEN_4 = _T_175 ? io_enable_bits_control : enable_R_control; // @[PhiNode.scala 222:26]
  assign _GEN_5 = _T_175 ? 1'h1 : enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_178 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_178 ? io_InData_0_bits_taskID : in_data_R_0_taskID; // @[PhiNode.scala 230:29]
  assign _GEN_8 = _T_178 ? 32'h0 : in_data_R_0_data; // @[PhiNode.scala 230:29]
  assign _GEN_9 = _T_178 ? 1'h1 : in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_181 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_181 ? io_InData_1_bits_taskID : in_data_R_1_taskID; // @[PhiNode.scala 230:29]
  assign _GEN_12 = _T_181 ? io_InData_1_bits_data : in_data_R_1_data; // @[PhiNode.scala 230:29]
  assign _GEN_13 = _T_181 ? 1'h1 : in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_183 = mask_R[0]; // @[Bitwise.scala 109:18]
  assign _T_184 = mask_R[1]; // @[Bitwise.scala 109:44]
  assign _T_185 = {_T_183,_T_184}; // @[Cat.scala 30:58]
  assign sel = _T_185[1]; // @[CircuitMath.scala 30:8]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[PhiNode.scala 250:43]
  assign _GEN_18 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 253:20]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_198 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_20 = _T_198 ? 1'h1 : fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_198 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_201 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_22 = _T_201 ? 1'h1 : fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_201 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_198; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_201; // @[PhiNode.scala 265:74]
  assign _T_207 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_208 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_209 = enable_valid_R & _T_208; // @[PhiNode.scala 277:27]
  assign _GEN_24 = enable_R_control ? 2'h1 : 2'h2; // @[PhiNode.scala 279:32]
  assign _GEN_25 = _T_209 ? 1'h1 : _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_26 = _T_209 ? 1'h1 : _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_27 = _T_209 ? _GEN_24 : state; // @[PhiNode.scala 277:46]
  assign _T_212 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_213 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _GEN_28 = _T_213 ? 32'h0 : _GEN_8; // @[PhiNode.scala 299:37]
  assign _GEN_29 = _T_213 ? 10'h0 : _GEN_7; // @[PhiNode.scala 299:37]
  assign _GEN_31 = _T_213 ? 32'h0 : _GEN_12; // @[PhiNode.scala 299:37]
  assign _GEN_32 = _T_213 ? 10'h0 : _GEN_11; // @[PhiNode.scala 299:37]
  assign _GEN_34 = _T_213 ? 1'h0 : _GEN_9; // @[PhiNode.scala 299:37]
  assign _GEN_35 = _T_213 ? 1'h0 : _GEN_13; // @[PhiNode.scala 299:37]
  assign _GEN_36 = _T_213 ? 2'h0 : _GEN_1; // @[PhiNode.scala 299:37]
  assign _GEN_37 = _T_213 ? 1'h0 : _GEN_2; // @[PhiNode.scala 299:37]
  assign _GEN_38 = _T_213 ? 1'h0 : _GEN_4; // @[PhiNode.scala 299:37]
  assign _GEN_39 = _T_213 ? 10'h0 : _GEN_3; // @[PhiNode.scala 299:37]
  assign _GEN_40 = _T_213 ? 1'h0 : _GEN_5; // @[PhiNode.scala 299:37]
  assign _GEN_41 = _T_213 ? 1'h0 : _GEN_20; // @[PhiNode.scala 299:37]
  assign _GEN_42 = _T_213 ? 1'h0 : _GEN_22; // @[PhiNode.scala 299:37]
  assign _GEN_43 = _T_213 ? 2'h0 : state; // @[PhiNode.scala 299:37]
  assign _T_235 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_60 = _T_235 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_64 = _T_235 ? task_input : _GEN_18; // @[Conditional.scala 39:67]
  assign _GEN_66 = _T_235 ? _GEN_28 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_67 = _T_235 ? _GEN_29 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_69 = _T_235 ? _GEN_31 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_70 = _T_235 ? _GEN_32 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_72 = _T_235 ? _GEN_34 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_73 = _T_235 ? _GEN_35 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_74 = _T_235 ? _GEN_36 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_75 = _T_235 ? _GEN_37 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_76 = _T_235 ? _GEN_38 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_77 = _T_235 ? _GEN_39 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_78 = _T_235 ? _GEN_40 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_79 = _T_235 ? _GEN_41 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_80 = _T_235 ? _GEN_42 : _GEN_22; // @[Conditional.scala 39:67]
  assign _GEN_81 = _T_235 ? _GEN_43 : state; // @[Conditional.scala 39:67]
  assign _GEN_82 = _T_212 ? _GEN_28 : _GEN_66; // @[Conditional.scala 39:67]
  assign _GEN_83 = _T_212 ? _GEN_29 : _GEN_67; // @[Conditional.scala 39:67]
  assign _GEN_85 = _T_212 ? _GEN_31 : _GEN_69; // @[Conditional.scala 39:67]
  assign _GEN_86 = _T_212 ? _GEN_32 : _GEN_70; // @[Conditional.scala 39:67]
  assign _GEN_88 = _T_212 ? _GEN_34 : _GEN_72; // @[Conditional.scala 39:67]
  assign _GEN_89 = _T_212 ? _GEN_35 : _GEN_73; // @[Conditional.scala 39:67]
  assign _GEN_90 = _T_212 ? _GEN_36 : _GEN_74; // @[Conditional.scala 39:67]
  assign _GEN_91 = _T_212 ? _GEN_37 : _GEN_75; // @[Conditional.scala 39:67]
  assign _GEN_92 = _T_212 ? _GEN_38 : _GEN_76; // @[Conditional.scala 39:67]
  assign _GEN_93 = _T_212 ? _GEN_39 : _GEN_77; // @[Conditional.scala 39:67]
  assign _GEN_94 = _T_212 ? _GEN_40 : _GEN_78; // @[Conditional.scala 39:67]
  assign _GEN_95 = _T_212 ? _GEN_41 : _GEN_79; // @[Conditional.scala 39:67]
  assign _GEN_96 = _T_212 ? _GEN_42 : _GEN_80; // @[Conditional.scala 39:67]
  assign _GEN_97 = _T_212 ? _GEN_43 : _GEN_81; // @[Conditional.scala 39:67]
  assign _GEN_98 = _T_212 ? _GEN_19 : _GEN_60; // @[Conditional.scala 39:67]
  assign _GEN_102 = _T_212 ? _GEN_18 : _GEN_64; // @[Conditional.scala 39:67]
  assign _GEN_104 = _T_207 ? _GEN_25 : _GEN_21; // @[Conditional.scala 40:58]
  assign _GEN_105 = _T_207 ? _GEN_26 : _GEN_23; // @[Conditional.scala 40:58]
  assign _GEN_106 = _T_207 ? _GEN_27 : _GEN_97; // @[Conditional.scala 40:58]
  assign _GEN_107 = _T_207 ? _GEN_8 : _GEN_82; // @[Conditional.scala 40:58]
  assign _GEN_108 = _T_207 ? _GEN_7 : _GEN_83; // @[Conditional.scala 40:58]
  assign _GEN_110 = _T_207 ? _GEN_12 : _GEN_85; // @[Conditional.scala 40:58]
  assign _GEN_111 = _T_207 ? _GEN_11 : _GEN_86; // @[Conditional.scala 40:58]
  assign _GEN_113 = _T_207 ? _GEN_9 : _GEN_88; // @[Conditional.scala 40:58]
  assign _GEN_114 = _T_207 ? _GEN_13 : _GEN_89; // @[Conditional.scala 40:58]
  assign _GEN_115 = _T_207 ? _GEN_1 : _GEN_90; // @[Conditional.scala 40:58]
  assign _GEN_116 = _T_207 ? _GEN_2 : _GEN_91; // @[Conditional.scala 40:58]
  assign _GEN_117 = _T_207 ? _GEN_4 : _GEN_92; // @[Conditional.scala 40:58]
  assign _GEN_118 = _T_207 ? _GEN_3 : _GEN_93; // @[Conditional.scala 40:58]
  assign _GEN_119 = _T_207 ? _GEN_5 : _GEN_94; // @[Conditional.scala 40:58]
  assign _GEN_120 = _T_207 ? _GEN_20 : _GEN_95; // @[Conditional.scala 40:58]
  assign _GEN_121 = _T_207 ? _GEN_22 : _GEN_96; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_207 ? _GEN_19 : _GEN_98; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_taskID = _T_207 ? _GEN_18 : _GEN_102; // @[PhiNode.scala 253:20 PhiNode.scala 326:44]
  assign io_Out_1_bits_data = _T_207 ? _GEN_19 : _GEN_98; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enable_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enable_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mask_R = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      in_data_R_0_taskID <= 10'h0;
    end else begin
      if (_T_207) begin
        if (_T_178) begin
          in_data_R_0_taskID <= io_InData_0_bits_taskID;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            in_data_R_0_taskID <= 10'h0;
          end else begin
            if (_T_178) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              in_data_R_0_taskID <= 10'h0;
            end else begin
              if (_T_178) begin
                in_data_R_0_taskID <= io_InData_0_bits_taskID;
              end
            end
          end else begin
            if (_T_178) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_207) begin
        if (_T_178) begin
          in_data_R_0_data <= 32'h0;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_178) begin
              in_data_R_0_data <= 32'h0;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_178) begin
                in_data_R_0_data <= 32'h0;
              end
            end
          end else begin
            if (_T_178) begin
              in_data_R_0_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 10'h0;
    end else begin
      if (_T_207) begin
        if (_T_181) begin
          in_data_R_1_taskID <= io_InData_1_bits_taskID;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            in_data_R_1_taskID <= 10'h0;
          end else begin
            if (_T_181) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              in_data_R_1_taskID <= 10'h0;
            end else begin
              if (_T_181) begin
                in_data_R_1_taskID <= io_InData_1_bits_taskID;
              end
            end
          end else begin
            if (_T_181) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_207) begin
        if (_T_181) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_181) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_181) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_181) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_178) begin
          in_data_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            if (_T_178) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              if (_T_178) begin
                in_data_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_178) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_181) begin
          in_data_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            if (_T_181) begin
              in_data_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              if (_T_181) begin
                in_data_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_181) begin
              in_data_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_207) begin
        if (_T_175) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_175) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_175) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_175) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_175) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_175) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_175) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_175) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_175) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_175) begin
              enable_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_175) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_175) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_207) begin
        if (_T_172) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_172) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_172) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_172) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_172) begin
          mask_valid_R <= 1'h1;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            mask_valid_R <= 1'h0;
          end else begin
            if (_T_172) begin
              mask_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              mask_valid_R <= 1'h0;
            end else begin
              if (_T_172) begin
                mask_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_172) begin
              mask_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_209) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_198) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_198) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_209) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_201) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_201) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_198) begin
          fire_R_0 <= 1'h1;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            fire_R_0 <= 1'h0;
          end else begin
            if (_T_198) begin
              fire_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              fire_R_0 <= 1'h0;
            end else begin
              if (_T_198) begin
                fire_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_198) begin
              fire_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_207) begin
        if (_T_201) begin
          fire_R_1 <= 1'h1;
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            fire_R_1 <= 1'h0;
          end else begin
            if (_T_201) begin
              fire_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              fire_R_1 <= 1'h0;
            end else begin
              if (_T_201) begin
                fire_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_201) begin
              fire_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_207) begin
        if (_T_209) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_212) begin
          if (_T_213) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_235) begin
            if (_T_213) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module UALU(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire [8:0] _T_21; // @[Alu.scala 108:45]
  wire [542:0] _GEN_0; // @[Alu.scala 108:36]
  wire [542:0] _T_22; // @[Alu.scala 108:36]
  assign _T_21 = io_in2[8:0]; // @[Alu.scala 108:45]
  assign _GEN_0 = {{511'd0}, io_in1}; // @[Alu.scala 108:36]
  assign _T_22 = _GEN_0 << _T_21; // @[Alu.scala 108:36]
  assign io_out = _T_22[31:0]; // @[Alu.scala 123:10]
endmodule
module ComputeNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? 32'h6 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h6;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UBranchNode_3(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_142; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_145; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_5;
  wire  _T_156; // @[Conditional.scala 37:30]
  wire  _GEN_6; // @[BranchNode.scala 611:46]
  wire  _GEN_7; // @[BranchNode.scala 611:46]
  wire  _T_168; // @[HandShaking.scala 656:24]
  wire  _T_170; // @[HandShaking.scala 656:24]
  wire  _T_171; // @[HandShaking.scala 656:50]
  wire  _T_173; // @[HandShaking.scala 656:50]
  wire  _T_174; // @[HandShaking.scala 656:29]
  wire  _GEN_8; // @[BranchNode.scala 631:26]
  wire  _GEN_9; // @[BranchNode.scala 631:26]
  wire  _GEN_10; // @[BranchNode.scala 631:26]
  wire  _GEN_11; // @[BranchNode.scala 631:26]
  wire [9:0] _GEN_12; // @[BranchNode.scala 631:26]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_21; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_23; // @[Conditional.scala 40:58]
  assign _T_142 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_142 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_142 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_145 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_145 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_145 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_145 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_156 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_6 = enable_valid_R ? 1'h1 : state; // @[BranchNode.scala 611:46]
  assign _GEN_7 = enable_valid_R ? 1'h1 : _GEN_1; // @[BranchNode.scala 611:46]
  assign _T_168 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_170 = _T_168 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_171 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_173 = _T_171 == 1'h0; // @[HandShaking.scala 656:50]
  assign _T_174 = _T_170 | _T_173; // @[HandShaking.scala 656:29]
  assign _GEN_8 = _T_174 ? 1'h0 : state; // @[BranchNode.scala 631:26]
  assign _GEN_9 = _T_174 ? 1'h0 : _GEN_0; // @[BranchNode.scala 631:26]
  assign _GEN_10 = _T_174 ? 1'h0 : _GEN_2; // @[BranchNode.scala 631:26]
  assign _GEN_11 = _T_174 ? 1'h0 : _GEN_3; // @[BranchNode.scala 631:26]
  assign _GEN_12 = _T_174 ? 10'h0 : _GEN_4; // @[BranchNode.scala 631:26]
  assign _GEN_13 = state ? _GEN_8 : state; // @[Conditional.scala 39:67]
  assign _GEN_14 = state ? _GEN_9 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_11 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_12 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_156 ? _GEN_6 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_156 ? _GEN_7 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_156 ? _GEN_0 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_156 ? _GEN_2 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_156 ? _GEN_3 : _GEN_16; // @[Conditional.scala 40:58]
  assign _GEN_23 = _T_156 ? _GEN_4 : _GEN_17; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 606:20]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 606:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_145) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_145) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_142) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_142) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_142) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_142) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_142) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module PhiFastNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [9:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [9:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [9:0]  io_Out_2_bits_taskID,
  output [31:0] io_Out_2_bits_data
);
  reg [9:0] in_data_R_0_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_0;
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [9:0] in_data_R_1_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_5;
  reg [9:0] enable_R_taskID; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_6;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_7;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_8;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_9;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_10;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_12;
  reg  out_valid_R_2; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_13;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_15;
  reg  fire_R_2; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_16;
  wire  _T_180; // @[Decoupled.scala 37:37]
  wire [1:0] _GEN_1; // @[PhiNode.scala 215:24]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_183; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[PhiNode.scala 222:26]
  wire  _GEN_4; // @[PhiNode.scala 222:26]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_186; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[PhiNode.scala 230:29]
  wire [31:0] _GEN_8; // @[PhiNode.scala 230:29]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_189; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[PhiNode.scala 230:29]
  wire [31:0] _GEN_12; // @[PhiNode.scala 230:29]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_191; // @[Bitwise.scala 109:18]
  wire  _T_192; // @[Bitwise.scala 109:44]
  wire [1:0] _T_193; // @[Cat.scala 30:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [9:0] task_input; // @[PhiNode.scala 250:43]
  wire [9:0] _GEN_18; // @[PhiNode.scala 253:20]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_209; // @[Decoupled.scala 37:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_212; // @[Decoupled.scala 37:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  _T_215; // @[Decoupled.scala 37:37]
  wire  _GEN_24; // @[PhiNode.scala 258:26]
  wire  _GEN_25; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  wire  fire_mask_2; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_17;
  wire  _T_222; // @[Conditional.scala 37:30]
  wire  _T_223; // @[PhiNode.scala 268:37]
  wire  _T_224; // @[PhiNode.scala 277:27]
  wire [1:0] _GEN_26; // @[PhiNode.scala 279:32]
  wire  _GEN_27; // @[PhiNode.scala 277:46]
  wire  _GEN_28; // @[PhiNode.scala 277:46]
  wire  _GEN_29; // @[PhiNode.scala 277:46]
  wire [1:0] _GEN_30; // @[PhiNode.scala 277:46]
  wire  _T_228; // @[Conditional.scala 37:30]
  wire  _T_229; // @[PhiNode.scala 299:31]
  wire  _T_230; // @[PhiNode.scala 299:31]
  wire [31:0] _GEN_31; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_32; // @[PhiNode.scala 299:37]
  wire [31:0] _GEN_34; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_35; // @[PhiNode.scala 299:37]
  wire  _GEN_37; // @[PhiNode.scala 299:37]
  wire  _GEN_38; // @[PhiNode.scala 299:37]
  wire [1:0] _GEN_39; // @[PhiNode.scala 299:37]
  wire  _GEN_40; // @[PhiNode.scala 299:37]
  wire  _GEN_41; // @[PhiNode.scala 299:37]
  wire [9:0] _GEN_42; // @[PhiNode.scala 299:37]
  wire  _GEN_43; // @[PhiNode.scala 299:37]
  wire  _GEN_44; // @[PhiNode.scala 299:37]
  wire  _GEN_45; // @[PhiNode.scala 299:37]
  wire  _GEN_46; // @[PhiNode.scala 299:37]
  wire [1:0] _GEN_47; // @[PhiNode.scala 299:37]
  wire  _T_253; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_65; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_71; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_74; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_75; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_77; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_78; // @[Conditional.scala 39:67]
  wire  _GEN_80; // @[Conditional.scala 39:67]
  wire  _GEN_81; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_82; // @[Conditional.scala 39:67]
  wire  _GEN_83; // @[Conditional.scala 39:67]
  wire  _GEN_84; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_85; // @[Conditional.scala 39:67]
  wire  _GEN_86; // @[Conditional.scala 39:67]
  wire  _GEN_87; // @[Conditional.scala 39:67]
  wire  _GEN_88; // @[Conditional.scala 39:67]
  wire  _GEN_89; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_90; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_91; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_92; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_94; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_97; // @[Conditional.scala 39:67]
  wire  _GEN_98; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_99; // @[Conditional.scala 39:67]
  wire  _GEN_100; // @[Conditional.scala 39:67]
  wire  _GEN_101; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_102; // @[Conditional.scala 39:67]
  wire  _GEN_103; // @[Conditional.scala 39:67]
  wire  _GEN_104; // @[Conditional.scala 39:67]
  wire  _GEN_105; // @[Conditional.scala 39:67]
  wire  _GEN_106; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_107; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_114; // @[Conditional.scala 39:67]
  wire  _GEN_117; // @[Conditional.scala 40:58]
  wire  _GEN_118; // @[Conditional.scala 40:58]
  wire  _GEN_119; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_120; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_121; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_122; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_124; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_125; // @[Conditional.scala 40:58]
  wire  _GEN_127; // @[Conditional.scala 40:58]
  wire  _GEN_128; // @[Conditional.scala 40:58]
  wire [1:0] _GEN_129; // @[Conditional.scala 40:58]
  wire  _GEN_130; // @[Conditional.scala 40:58]
  wire  _GEN_131; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_132; // @[Conditional.scala 40:58]
  wire  _GEN_133; // @[Conditional.scala 40:58]
  wire  _GEN_134; // @[Conditional.scala 40:58]
  wire  _GEN_135; // @[Conditional.scala 40:58]
  wire  _GEN_136; // @[Conditional.scala 40:58]
  assign _T_180 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_180 ? io_Mask_bits : mask_R; // @[PhiNode.scala 215:24]
  assign _GEN_2 = _T_180 ? 1'h1 : mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_183 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_183 ? io_enable_bits_taskID : enable_R_taskID; // @[PhiNode.scala 222:26]
  assign _GEN_4 = _T_183 ? io_enable_bits_control : enable_R_control; // @[PhiNode.scala 222:26]
  assign _GEN_5 = _T_183 ? 1'h1 : enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_186 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_186 ? io_InData_0_bits_taskID : in_data_R_0_taskID; // @[PhiNode.scala 230:29]
  assign _GEN_8 = _T_186 ? 32'h0 : in_data_R_0_data; // @[PhiNode.scala 230:29]
  assign _GEN_9 = _T_186 ? 1'h1 : in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_189 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_189 ? io_InData_1_bits_taskID : in_data_R_1_taskID; // @[PhiNode.scala 230:29]
  assign _GEN_12 = _T_189 ? io_InData_1_bits_data : in_data_R_1_data; // @[PhiNode.scala 230:29]
  assign _GEN_13 = _T_189 ? 1'h1 : in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_191 = mask_R[0]; // @[Bitwise.scala 109:18]
  assign _T_192 = mask_R[1]; // @[Bitwise.scala 109:44]
  assign _T_193 = {_T_191,_T_192}; // @[Cat.scala 30:58]
  assign sel = _T_193[1]; // @[CircuitMath.scala 30:8]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[PhiNode.scala 250:43]
  assign _GEN_18 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 253:20]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_209 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_20 = _T_209 ? 1'h1 : fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_209 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_212 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_22 = _T_212 ? 1'h1 : fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_212 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign _T_215 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 37:37]
  assign _GEN_24 = _T_215 ? 1'h1 : fire_R_2; // @[PhiNode.scala 258:26]
  assign _GEN_25 = _T_215 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_209; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_212; // @[PhiNode.scala 265:74]
  assign fire_mask_2 = fire_R_2 | _T_215; // @[PhiNode.scala 265:74]
  assign _T_222 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_223 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_224 = enable_valid_R & _T_223; // @[PhiNode.scala 277:27]
  assign _GEN_26 = enable_R_control ? 2'h1 : 2'h2; // @[PhiNode.scala 279:32]
  assign _GEN_27 = _T_224 ? 1'h1 : _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_28 = _T_224 ? 1'h1 : _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_29 = _T_224 ? 1'h1 : _GEN_25; // @[PhiNode.scala 277:46]
  assign _GEN_30 = _T_224 ? _GEN_26 : state; // @[PhiNode.scala 277:46]
  assign _T_228 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_229 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_230 = _T_229 & fire_mask_2; // @[PhiNode.scala 299:31]
  assign _GEN_31 = _T_230 ? 32'h0 : _GEN_8; // @[PhiNode.scala 299:37]
  assign _GEN_32 = _T_230 ? 10'h0 : _GEN_7; // @[PhiNode.scala 299:37]
  assign _GEN_34 = _T_230 ? 32'h0 : _GEN_12; // @[PhiNode.scala 299:37]
  assign _GEN_35 = _T_230 ? 10'h0 : _GEN_11; // @[PhiNode.scala 299:37]
  assign _GEN_37 = _T_230 ? 1'h0 : _GEN_9; // @[PhiNode.scala 299:37]
  assign _GEN_38 = _T_230 ? 1'h0 : _GEN_13; // @[PhiNode.scala 299:37]
  assign _GEN_39 = _T_230 ? 2'h0 : _GEN_1; // @[PhiNode.scala 299:37]
  assign _GEN_40 = _T_230 ? 1'h0 : _GEN_2; // @[PhiNode.scala 299:37]
  assign _GEN_41 = _T_230 ? 1'h0 : _GEN_4; // @[PhiNode.scala 299:37]
  assign _GEN_42 = _T_230 ? 10'h0 : _GEN_3; // @[PhiNode.scala 299:37]
  assign _GEN_43 = _T_230 ? 1'h0 : _GEN_5; // @[PhiNode.scala 299:37]
  assign _GEN_44 = _T_230 ? 1'h0 : _GEN_20; // @[PhiNode.scala 299:37]
  assign _GEN_45 = _T_230 ? 1'h0 : _GEN_22; // @[PhiNode.scala 299:37]
  assign _GEN_46 = _T_230 ? 1'h0 : _GEN_24; // @[PhiNode.scala 299:37]
  assign _GEN_47 = _T_230 ? 2'h0 : state; // @[PhiNode.scala 299:37]
  assign _T_253 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_65 = _T_253 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_71 = _T_253 ? task_input : _GEN_18; // @[Conditional.scala 39:67]
  assign _GEN_74 = _T_253 ? _GEN_31 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_75 = _T_253 ? _GEN_32 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_77 = _T_253 ? _GEN_34 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_78 = _T_253 ? _GEN_35 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_80 = _T_253 ? _GEN_37 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_81 = _T_253 ? _GEN_38 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_82 = _T_253 ? _GEN_39 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_83 = _T_253 ? _GEN_40 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_84 = _T_253 ? _GEN_41 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_85 = _T_253 ? _GEN_42 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_86 = _T_253 ? _GEN_43 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_87 = _T_253 ? _GEN_44 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_88 = _T_253 ? _GEN_45 : _GEN_22; // @[Conditional.scala 39:67]
  assign _GEN_89 = _T_253 ? _GEN_46 : _GEN_24; // @[Conditional.scala 39:67]
  assign _GEN_90 = _T_253 ? _GEN_47 : state; // @[Conditional.scala 39:67]
  assign _GEN_91 = _T_228 ? _GEN_31 : _GEN_74; // @[Conditional.scala 39:67]
  assign _GEN_92 = _T_228 ? _GEN_32 : _GEN_75; // @[Conditional.scala 39:67]
  assign _GEN_94 = _T_228 ? _GEN_34 : _GEN_77; // @[Conditional.scala 39:67]
  assign _GEN_95 = _T_228 ? _GEN_35 : _GEN_78; // @[Conditional.scala 39:67]
  assign _GEN_97 = _T_228 ? _GEN_37 : _GEN_80; // @[Conditional.scala 39:67]
  assign _GEN_98 = _T_228 ? _GEN_38 : _GEN_81; // @[Conditional.scala 39:67]
  assign _GEN_99 = _T_228 ? _GEN_39 : _GEN_82; // @[Conditional.scala 39:67]
  assign _GEN_100 = _T_228 ? _GEN_40 : _GEN_83; // @[Conditional.scala 39:67]
  assign _GEN_101 = _T_228 ? _GEN_41 : _GEN_84; // @[Conditional.scala 39:67]
  assign _GEN_102 = _T_228 ? _GEN_42 : _GEN_85; // @[Conditional.scala 39:67]
  assign _GEN_103 = _T_228 ? _GEN_43 : _GEN_86; // @[Conditional.scala 39:67]
  assign _GEN_104 = _T_228 ? _GEN_44 : _GEN_87; // @[Conditional.scala 39:67]
  assign _GEN_105 = _T_228 ? _GEN_45 : _GEN_88; // @[Conditional.scala 39:67]
  assign _GEN_106 = _T_228 ? _GEN_46 : _GEN_89; // @[Conditional.scala 39:67]
  assign _GEN_107 = _T_228 ? _GEN_47 : _GEN_90; // @[Conditional.scala 39:67]
  assign _GEN_108 = _T_228 ? _GEN_19 : _GEN_65; // @[Conditional.scala 39:67]
  assign _GEN_114 = _T_228 ? _GEN_18 : _GEN_71; // @[Conditional.scala 39:67]
  assign _GEN_117 = _T_222 ? _GEN_27 : _GEN_21; // @[Conditional.scala 40:58]
  assign _GEN_118 = _T_222 ? _GEN_28 : _GEN_23; // @[Conditional.scala 40:58]
  assign _GEN_119 = _T_222 ? _GEN_29 : _GEN_25; // @[Conditional.scala 40:58]
  assign _GEN_120 = _T_222 ? _GEN_30 : _GEN_107; // @[Conditional.scala 40:58]
  assign _GEN_121 = _T_222 ? _GEN_8 : _GEN_91; // @[Conditional.scala 40:58]
  assign _GEN_122 = _T_222 ? _GEN_7 : _GEN_92; // @[Conditional.scala 40:58]
  assign _GEN_124 = _T_222 ? _GEN_12 : _GEN_94; // @[Conditional.scala 40:58]
  assign _GEN_125 = _T_222 ? _GEN_11 : _GEN_95; // @[Conditional.scala 40:58]
  assign _GEN_127 = _T_222 ? _GEN_9 : _GEN_97; // @[Conditional.scala 40:58]
  assign _GEN_128 = _T_222 ? _GEN_13 : _GEN_98; // @[Conditional.scala 40:58]
  assign _GEN_129 = _T_222 ? _GEN_1 : _GEN_99; // @[Conditional.scala 40:58]
  assign _GEN_130 = _T_222 ? _GEN_2 : _GEN_100; // @[Conditional.scala 40:58]
  assign _GEN_131 = _T_222 ? _GEN_4 : _GEN_101; // @[Conditional.scala 40:58]
  assign _GEN_132 = _T_222 ? _GEN_3 : _GEN_102; // @[Conditional.scala 40:58]
  assign _GEN_133 = _T_222 ? _GEN_5 : _GEN_103; // @[Conditional.scala 40:58]
  assign _GEN_134 = _T_222 ? _GEN_20 : _GEN_104; // @[Conditional.scala 40:58]
  assign _GEN_135 = _T_222 ? _GEN_22 : _GEN_105; // @[Conditional.scala 40:58]
  assign _GEN_136 = _T_222 ? _GEN_24 : _GEN_106; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_222 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_222 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 254:21]
  assign io_Out_2_bits_taskID = _T_222 ? _GEN_18 : _GEN_114; // @[PhiNode.scala 253:20 PhiNode.scala 326:44]
  assign io_Out_2_bits_data = _T_222 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 324:42]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enable_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enable_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mask_R = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fire_R_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  fire_R_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  state = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      in_data_R_0_taskID <= 10'h0;
    end else begin
      if (_T_222) begin
        if (_T_186) begin
          in_data_R_0_taskID <= io_InData_0_bits_taskID;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            in_data_R_0_taskID <= 10'h0;
          end else begin
            if (_T_186) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              in_data_R_0_taskID <= 10'h0;
            end else begin
              if (_T_186) begin
                in_data_R_0_taskID <= io_InData_0_bits_taskID;
              end
            end
          end else begin
            if (_T_186) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_222) begin
        if (_T_186) begin
          in_data_R_0_data <= 32'h0;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_186) begin
              in_data_R_0_data <= 32'h0;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_186) begin
                in_data_R_0_data <= 32'h0;
              end
            end
          end else begin
            if (_T_186) begin
              in_data_R_0_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 10'h0;
    end else begin
      if (_T_222) begin
        if (_T_189) begin
          in_data_R_1_taskID <= io_InData_1_bits_taskID;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            in_data_R_1_taskID <= 10'h0;
          end else begin
            if (_T_189) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              in_data_R_1_taskID <= 10'h0;
            end else begin
              if (_T_189) begin
                in_data_R_1_taskID <= io_InData_1_bits_taskID;
              end
            end
          end else begin
            if (_T_189) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_222) begin
        if (_T_189) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_189) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_189) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_189) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_186) begin
          in_data_valid_R_0 <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            if (_T_186) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              if (_T_186) begin
                in_data_valid_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_186) begin
              in_data_valid_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_189) begin
          in_data_valid_R_1 <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            if (_T_189) begin
              in_data_valid_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              if (_T_189) begin
                in_data_valid_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_189) begin
              in_data_valid_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_222) begin
        if (_T_183) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_183) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              enable_R_taskID <= 10'h0;
            end else begin
              if (_T_183) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_183) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_183) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_183) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_183) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_183) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_183) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_183) begin
              enable_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_183) begin
                enable_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_183) begin
              enable_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_222) begin
        if (_T_180) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_180) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_180) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_180) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_180) begin
          mask_valid_R <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            mask_valid_R <= 1'h0;
          end else begin
            if (_T_180) begin
              mask_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              mask_valid_R <= 1'h0;
            end else begin
              if (_T_180) begin
                mask_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_180) begin
              mask_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_224) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_209) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_209) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_224) begin
          out_valid_R_1 <= 1'h1;
        end else begin
          if (_T_212) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_212) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_224) begin
          out_valid_R_2 <= 1'h1;
        end else begin
          if (_T_215) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_215) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_209) begin
          fire_R_0 <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            fire_R_0 <= 1'h0;
          end else begin
            if (_T_209) begin
              fire_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              fire_R_0 <= 1'h0;
            end else begin
              if (_T_209) begin
                fire_R_0 <= 1'h1;
              end
            end
          end else begin
            if (_T_209) begin
              fire_R_0 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_212) begin
          fire_R_1 <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            fire_R_1 <= 1'h0;
          end else begin
            if (_T_212) begin
              fire_R_1 <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              fire_R_1 <= 1'h0;
            end else begin
              if (_T_212) begin
                fire_R_1 <= 1'h1;
              end
            end
          end else begin
            if (_T_212) begin
              fire_R_1 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else begin
      if (_T_222) begin
        if (_T_215) begin
          fire_R_2 <= 1'h1;
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            fire_R_2 <= 1'h0;
          end else begin
            if (_T_215) begin
              fire_R_2 <= 1'h1;
            end
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              fire_R_2 <= 1'h0;
            end else begin
              if (_T_215) begin
                fire_R_2 <= 1'h1;
              end
            end
          end else begin
            if (_T_215) begin
              fire_R_2 <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_222) begin
        if (_T_224) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_228) begin
          if (_T_230) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_253) begin
            if (_T_230) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module UALU_1(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire [32:0] _T_11; // @[Alu.scala 102:30]
  assign _T_11 = io_in1 + io_in2; // @[Alu.scala 102:30]
  assign io_out = io_in1 + io_in2; // @[Alu.scala 123:10]
endmodule
module ComputeNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? 32'h6 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h6;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module GepNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [9:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] base_addr_R_taskID; // @[GepNode.scala 892:28]
  reg [31:0] _RAND_4;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 892:28]
  reg [31:0] _RAND_5;
  reg  base_addr_valid_R; // @[GepNode.scala 893:34]
  reg [31:0] _RAND_6;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 896:39]
  reg [31:0] _RAND_7;
  reg  idx_valid_R_0; // @[GepNode.scala 897:45]
  reg [31:0] _RAND_8;
  reg  state; // @[GepNode.scala 901:22]
  reg [31:0] _RAND_9;
  wire  _T_119; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[GepNode.scala 917:31]
  wire [31:0] _GEN_8; // @[GepNode.scala 917:31]
  wire  _GEN_9; // @[GepNode.scala 917:31]
  wire  _T_122; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[GepNode.scala 924:28]
  wire  _GEN_13; // @[GepNode.scala 924:28]
  wire [35:0] seek_value; // @[GepNode.scala 932:21]
  wire [35:0] _GEN_54; // @[GepNode.scala 940:35]
  wire [36:0] _T_125; // @[GepNode.scala 940:35]
  wire [35:0] data_out; // @[GepNode.scala 940:35]
  wire  _T_126; // @[Conditional.scala 37:30]
  wire  _T_127; // @[GepNode.scala 958:42]
  wire  _GEN_14; // @[GepNode.scala 958:64]
  wire  _GEN_15; // @[GepNode.scala 958:64]
  wire  _GEN_16; // @[GepNode.scala 957:32]
  wire  _GEN_17; // @[GepNode.scala 957:32]
  wire  _GEN_18; // @[GepNode.scala 956:28]
  wire  _GEN_19; // @[GepNode.scala 956:28]
  wire  _T_132; // @[HandShaking.scala 222:83]
  wire [31:0] _GEN_20; // @[GepNode.scala 970:26]
  wire [31:0] _GEN_23; // @[GepNode.scala 970:26]
  wire [9:0] _GEN_24; // @[GepNode.scala 970:26]
  wire  _GEN_26; // @[GepNode.scala 970:26]
  wire  _GEN_27; // @[GepNode.scala 970:26]
  wire  _GEN_28; // @[GepNode.scala 970:26]
  wire  _GEN_29; // @[GepNode.scala 970:26]
  wire  _GEN_30; // @[GepNode.scala 970:26]
  wire [31:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_34; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_44; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_47; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  assign _T_88 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_88 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_88 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_119 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_119 ? io_baseAddress_bits_taskID : base_addr_R_taskID; // @[GepNode.scala 917:31]
  assign _GEN_8 = _T_119 ? io_baseAddress_bits_data : base_addr_R_data; // @[GepNode.scala 917:31]
  assign _GEN_9 = _T_119 ? 1'h1 : base_addr_valid_R; // @[GepNode.scala 917:31]
  assign _T_122 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_122 ? io_idx_0_bits_data : idx_R_0_data; // @[GepNode.scala 924:28]
  assign _GEN_13 = _T_122 ? 1'h1 : idx_valid_R_0; // @[GepNode.scala 924:28]
  assign seek_value = idx_R_0_data * 32'h8; // @[GepNode.scala 932:21]
  assign _GEN_54 = {{4'd0}, base_addr_R_data}; // @[GepNode.scala 940:35]
  assign _T_125 = _GEN_54 + seek_value; // @[GepNode.scala 940:35]
  assign data_out = _GEN_54 + seek_value; // @[GepNode.scala 940:35]
  assign _T_126 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_127 = idx_valid_R_0 & base_addr_valid_R; // @[GepNode.scala 958:42]
  assign _GEN_14 = _T_127 ? 1'h1 : _GEN_1; // @[GepNode.scala 958:64]
  assign _GEN_15 = _T_127 ? 1'h1 : state; // @[GepNode.scala 958:64]
  assign _GEN_16 = enable_R_control ? _GEN_14 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_17 = enable_R_control ? _GEN_15 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_18 = enable_valid_R ? _GEN_16 : _GEN_1; // @[GepNode.scala 956:28]
  assign _GEN_19 = enable_valid_R ? _GEN_17 : state; // @[GepNode.scala 956:28]
  assign _T_132 = out_ready_R_0 | _T_88; // @[HandShaking.scala 222:83]
  assign _GEN_20 = _T_132 ? 32'h0 : _GEN_12; // @[GepNode.scala 970:26]
  assign _GEN_23 = _T_132 ? 32'h0 : _GEN_8; // @[GepNode.scala 970:26]
  assign _GEN_24 = _T_132 ? 10'h0 : _GEN_7; // @[GepNode.scala 970:26]
  assign _GEN_26 = _T_132 ? 1'h0 : _GEN_13; // @[GepNode.scala 970:26]
  assign _GEN_27 = _T_132 ? 1'h0 : _GEN_9; // @[GepNode.scala 970:26]
  assign _GEN_28 = _T_132 ? 1'h0 : state; // @[GepNode.scala 970:26]
  assign _GEN_29 = _T_132 ? 1'h0 : _GEN_0; // @[GepNode.scala 970:26]
  assign _GEN_30 = _T_132 ? 1'h0 : _GEN_2; // @[GepNode.scala 970:26]
  assign _GEN_31 = state ? _GEN_20 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_23 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_24 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_26 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_28 : state; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_29 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_41 = state ? _GEN_30 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_126 ? _GEN_18 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_126 ? _GEN_19 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_126 ? _GEN_12 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_126 ? _GEN_8 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_126 ? _GEN_7 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_126 ? _GEN_13 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_126 ? _GEN_9 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_126 ? _GEN_0 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_126 ? _GEN_2 : _GEN_41; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 945:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 946:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 944:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 916:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 923:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  base_addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  idx_R_0_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_88) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_126) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_127) begin
              out_valid_R_0 <= 1'h1;
            end else begin
              if (_T_88) begin
                out_valid_R_0 <= 1'h0;
              end
            end
          end else begin
            out_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_88) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      base_addr_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        if (_T_119) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            base_addr_R_taskID <= 10'h0;
          end else begin
            if (_T_119) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_119) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_119) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_119) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_119) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_119) begin
          base_addr_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            if (_T_119) begin
              base_addr_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_119) begin
            base_addr_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_122) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_122) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_122) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_122) begin
          idx_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            if (_T_122) begin
              idx_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_122) begin
            idx_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_126) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_127) begin
              state <= 1'h1;
            end
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UnTypLoad(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [9:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [9:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_165; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_168; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_5;
  reg [9:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_8;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_10;
  wire  _T_196; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_6; // @[LoadSimple.scala 81:27]
  wire [9:0] _GEN_7; // @[LoadSimple.scala 81:27]
  wire  _GEN_8; // @[LoadSimple.scala 81:27]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  _T_199; // @[HandShaking.scala 656:24]
  wire  _T_201; // @[HandShaking.scala 656:24]
  wire  _T_202; // @[HandShaking.scala 656:50]
  wire  _T_204; // @[HandShaking.scala 656:50]
  wire  complete; // @[HandShaking.scala 656:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_211; // @[Conditional.scala 37:30]
  wire  _T_212; // @[LoadSimple.scala 119:27]
  wire  _T_213; // @[LoadSimple.scala 120:31]
  wire [1:0] _GEN_10; // @[LoadSimple.scala 122:33]
  wire [1:0] _GEN_12; // @[LoadSimple.scala 120:45]
  wire  _GEN_14; // @[LoadSimple.scala 120:45]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire [1:0] _GEN_16; // @[LoadSimple.scala 119:44]
  wire  _GEN_18; // @[LoadSimple.scala 119:44]
  wire  _T_224; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_19; // @[LoadSimple.scala 135:30]
  wire  _GEN_21; // @[LoadSimple.scala 135:30]
  wire [1:0] _GEN_22; // @[LoadSimple.scala 135:30]
  wire  _T_234; // @[Conditional.scala 37:30]
  wire  _GEN_23; // @[LoadSimple.scala 149:22]
  wire  _GEN_25; // @[LoadSimple.scala 149:22]
  wire  _GEN_26; // @[LoadSimple.scala 149:22]
  wire [1:0] _GEN_27; // @[LoadSimple.scala 149:22]
  wire  _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  assign _T_165 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_165 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_165 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_168 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_168 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_168 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_168 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_196 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_196 ? io_GepAddr_bits_data : addr_R_data; // @[LoadSimple.scala 81:27]
  assign _GEN_7 = _T_196 ? io_GepAddr_bits_taskID : addr_R_taskID; // @[LoadSimple.scala 81:27]
  assign _GEN_8 = _T_196 ? io_GepAddr_bits_predicate : addr_R_predicate; // @[LoadSimple.scala 81:27]
  assign _GEN_9 = _T_196 ? 1'h1 : addr_valid_R; // @[LoadSimple.scala 81:27]
  assign _T_199 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_201 = _T_199 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_202 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_204 = _T_202 == 1'h0; // @[HandShaking.scala 656:50]
  assign complete = _T_201 | _T_204; // @[HandShaking.scala 656:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_211 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_212 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_213 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _GEN_10 = io_memReq_ready ? 2'h1 : state; // @[LoadSimple.scala 122:33]
  assign _GEN_12 = _T_213 ? _GEN_10 : 2'h2; // @[LoadSimple.scala 120:45]
  assign _GEN_14 = _T_213 ? _GEN_1 : 1'h1; // @[LoadSimple.scala 120:45]
  assign _GEN_15 = _T_212 ? _T_213 : 1'h0; // @[LoadSimple.scala 119:44]
  assign _GEN_16 = _T_212 ? _GEN_12 : state; // @[LoadSimple.scala 119:44]
  assign _GEN_18 = _T_212 ? _GEN_14 : _GEN_1; // @[LoadSimple.scala 119:44]
  assign _T_224 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _GEN_19 = io_memResp_valid ? io_memResp_data : data_R_data; // @[LoadSimple.scala 135:30]
  assign _GEN_21 = io_memResp_valid ? 1'h1 : _GEN_1; // @[LoadSimple.scala 135:30]
  assign _GEN_22 = io_memResp_valid ? 2'h2 : state; // @[LoadSimple.scala 135:30]
  assign _T_234 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_23 = complete ? 1'h0 : _GEN_9; // @[LoadSimple.scala 149:22]
  assign _GEN_25 = complete ? 1'h0 : _GEN_0; // @[LoadSimple.scala 149:22]
  assign _GEN_26 = complete ? 1'h0 : _GEN_2; // @[LoadSimple.scala 149:22]
  assign _GEN_27 = complete ? 2'h0 : state; // @[LoadSimple.scala 149:22]
  assign _GEN_28 = _T_234 ? _GEN_23 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_234 ? _GEN_25 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_234 ? _GEN_26 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_234 ? _GEN_27 : state; // @[Conditional.scala 39:67]
  assign _GEN_33 = _T_224 ? _GEN_19 : data_R_data; // @[Conditional.scala 39:67]
  assign _GEN_35 = _T_224 ? _GEN_21 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_224 ? _GEN_22 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_224 ? _GEN_9 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_224 ? _GEN_0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_40 = _T_224 ? _GEN_2 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_211 ? _GEN_16 : _GEN_36; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_211 ? _GEN_18 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_211 ? data_R_data : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_211 ? _GEN_9 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_211 ? _GEN_0 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_211 ? _GEN_2 : _GEN_40; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = addr_R_taskID | enable_R_taskID; // @[LoadSimple.scala 97:20 LoadSimple.scala 99:27]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_211 ? _GEN_15 : 1'h0; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_predicate = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_168) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_168) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_168) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_224) begin
          if (_T_168) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_168) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_168) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_165) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_224) begin
          if (_T_165) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_165) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_165) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_212) begin
          if (_T_213) begin
            if (_T_165) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_165) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_165) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_165) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_196) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 10'h0;
    end else begin
      if (_T_196) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_196) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_196) begin
          addr_valid_R <= 1'h1;
        end
      end else begin
        if (_T_224) begin
          if (_T_196) begin
            addr_valid_R <= 1'h1;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              if (_T_196) begin
                addr_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_196) begin
              addr_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_211)) begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_211) begin
        if (_T_212) begin
          if (_T_213) begin
            if (io_memReq_ready) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module UBranchNode_4(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [9:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_142; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_145; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_5;
  wire  _T_156; // @[Conditional.scala 37:30]
  wire  _GEN_6; // @[BranchNode.scala 611:46]
  wire  _GEN_7; // @[BranchNode.scala 611:46]
  wire  _T_168; // @[HandShaking.scala 656:24]
  wire  _T_170; // @[HandShaking.scala 656:24]
  wire  _T_171; // @[HandShaking.scala 656:50]
  wire  _T_173; // @[HandShaking.scala 656:50]
  wire  _T_174; // @[HandShaking.scala 656:29]
  wire  _GEN_8; // @[BranchNode.scala 631:26]
  wire  _GEN_9; // @[BranchNode.scala 631:26]
  wire  _GEN_10; // @[BranchNode.scala 631:26]
  wire  _GEN_11; // @[BranchNode.scala 631:26]
  wire [9:0] _GEN_12; // @[BranchNode.scala 631:26]
  wire  _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_21; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_23; // @[Conditional.scala 40:58]
  assign _T_142 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_142 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_142 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_145 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_145 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_145 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_145 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_156 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_6 = enable_valid_R ? 1'h1 : state; // @[BranchNode.scala 611:46]
  assign _GEN_7 = enable_valid_R ? 1'h1 : _GEN_1; // @[BranchNode.scala 611:46]
  assign _T_168 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_170 = _T_168 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_171 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_173 = _T_171 == 1'h0; // @[HandShaking.scala 656:50]
  assign _T_174 = _T_170 | _T_173; // @[HandShaking.scala 656:29]
  assign _GEN_8 = _T_174 ? 1'h0 : state; // @[BranchNode.scala 631:26]
  assign _GEN_9 = _T_174 ? 1'h0 : _GEN_0; // @[BranchNode.scala 631:26]
  assign _GEN_10 = _T_174 ? 1'h0 : _GEN_2; // @[BranchNode.scala 631:26]
  assign _GEN_11 = _T_174 ? 1'h0 : _GEN_3; // @[BranchNode.scala 631:26]
  assign _GEN_12 = _T_174 ? 10'h0 : _GEN_4; // @[BranchNode.scala 631:26]
  assign _GEN_13 = state ? _GEN_8 : state; // @[Conditional.scala 39:67]
  assign _GEN_14 = state ? _GEN_9 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_11 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_12 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_156 ? _GEN_6 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_156 ? _GEN_7 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_156 ? _GEN_0 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_156 ? _GEN_2 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_156 ? _GEN_3 : _GEN_16; // @[Conditional.scala 40:58]
  assign _GEN_23 = _T_156 ? _GEN_4 : _GEN_17; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 606:20]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 606:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_145) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_145) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_145) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_145) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_145) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (_T_142) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_142) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_142) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= 1'h1;
        end else begin
          if (_T_142) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_142) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_156) begin
        if (enable_valid_R) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_174) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module GepNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [9:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] base_addr_R_taskID; // @[GepNode.scala 892:28]
  reg [31:0] _RAND_4;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 892:28]
  reg [31:0] _RAND_5;
  reg  base_addr_valid_R; // @[GepNode.scala 893:34]
  reg [31:0] _RAND_6;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 896:39]
  reg [31:0] _RAND_7;
  reg  idx_valid_R_0; // @[GepNode.scala 897:45]
  reg [31:0] _RAND_8;
  reg  state; // @[GepNode.scala 901:22]
  reg [31:0] _RAND_9;
  wire  _T_119; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[GepNode.scala 917:31]
  wire [31:0] _GEN_8; // @[GepNode.scala 917:31]
  wire  _GEN_9; // @[GepNode.scala 917:31]
  wire  _T_122; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[GepNode.scala 924:28]
  wire  _GEN_13; // @[GepNode.scala 924:28]
  wire [35:0] seek_value; // @[GepNode.scala 932:21]
  wire [35:0] _GEN_54; // @[GepNode.scala 940:35]
  wire [36:0] _T_125; // @[GepNode.scala 940:35]
  wire [35:0] data_out; // @[GepNode.scala 940:35]
  wire  _T_126; // @[Conditional.scala 37:30]
  wire  _T_127; // @[GepNode.scala 958:42]
  wire  _GEN_14; // @[GepNode.scala 958:64]
  wire  _GEN_15; // @[GepNode.scala 958:64]
  wire  _GEN_16; // @[GepNode.scala 957:32]
  wire  _GEN_17; // @[GepNode.scala 957:32]
  wire  _GEN_18; // @[GepNode.scala 956:28]
  wire  _GEN_19; // @[GepNode.scala 956:28]
  wire  _T_132; // @[HandShaking.scala 222:83]
  wire [31:0] _GEN_20; // @[GepNode.scala 970:26]
  wire [31:0] _GEN_23; // @[GepNode.scala 970:26]
  wire [9:0] _GEN_24; // @[GepNode.scala 970:26]
  wire  _GEN_26; // @[GepNode.scala 970:26]
  wire  _GEN_27; // @[GepNode.scala 970:26]
  wire  _GEN_28; // @[GepNode.scala 970:26]
  wire  _GEN_29; // @[GepNode.scala 970:26]
  wire  _GEN_30; // @[GepNode.scala 970:26]
  wire [31:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_34; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_44; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_47; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  assign _T_88 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_88 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_88 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_119 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_119 ? io_baseAddress_bits_taskID : base_addr_R_taskID; // @[GepNode.scala 917:31]
  assign _GEN_8 = _T_119 ? io_baseAddress_bits_data : base_addr_R_data; // @[GepNode.scala 917:31]
  assign _GEN_9 = _T_119 ? 1'h1 : base_addr_valid_R; // @[GepNode.scala 917:31]
  assign _T_122 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_122 ? io_idx_0_bits_data : idx_R_0_data; // @[GepNode.scala 924:28]
  assign _GEN_13 = _T_122 ? 1'h1 : idx_valid_R_0; // @[GepNode.scala 924:28]
  assign seek_value = idx_R_0_data * 32'h8; // @[GepNode.scala 932:21]
  assign _GEN_54 = {{4'd0}, base_addr_R_data}; // @[GepNode.scala 940:35]
  assign _T_125 = _GEN_54 + seek_value; // @[GepNode.scala 940:35]
  assign data_out = _GEN_54 + seek_value; // @[GepNode.scala 940:35]
  assign _T_126 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_127 = idx_valid_R_0 & base_addr_valid_R; // @[GepNode.scala 958:42]
  assign _GEN_14 = _T_127 ? 1'h1 : _GEN_1; // @[GepNode.scala 958:64]
  assign _GEN_15 = _T_127 ? 1'h1 : state; // @[GepNode.scala 958:64]
  assign _GEN_16 = enable_R_control ? _GEN_14 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_17 = enable_R_control ? _GEN_15 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_18 = enable_valid_R ? _GEN_16 : _GEN_1; // @[GepNode.scala 956:28]
  assign _GEN_19 = enable_valid_R ? _GEN_17 : state; // @[GepNode.scala 956:28]
  assign _T_132 = out_ready_R_0 | _T_88; // @[HandShaking.scala 222:83]
  assign _GEN_20 = _T_132 ? 32'h0 : _GEN_12; // @[GepNode.scala 970:26]
  assign _GEN_23 = _T_132 ? 32'h0 : _GEN_8; // @[GepNode.scala 970:26]
  assign _GEN_24 = _T_132 ? 10'h0 : _GEN_7; // @[GepNode.scala 970:26]
  assign _GEN_26 = _T_132 ? 1'h0 : _GEN_13; // @[GepNode.scala 970:26]
  assign _GEN_27 = _T_132 ? 1'h0 : _GEN_9; // @[GepNode.scala 970:26]
  assign _GEN_28 = _T_132 ? 1'h0 : state; // @[GepNode.scala 970:26]
  assign _GEN_29 = _T_132 ? 1'h0 : _GEN_0; // @[GepNode.scala 970:26]
  assign _GEN_30 = _T_132 ? 1'h0 : _GEN_2; // @[GepNode.scala 970:26]
  assign _GEN_31 = state ? _GEN_20 : _GEN_12; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_23 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_24 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_26 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_28 : state; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_29 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_41 = state ? _GEN_30 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_126 ? _GEN_18 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_126 ? _GEN_19 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_126 ? _GEN_12 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_126 ? _GEN_8 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_126 ? _GEN_7 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_126 ? _GEN_13 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_126 ? _GEN_9 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_126 ? _GEN_0 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_126 ? _GEN_2 : _GEN_41; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 945:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 946:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 944:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 916:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 923:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  base_addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  idx_R_0_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_88) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_126) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_127) begin
              out_valid_R_0 <= 1'h1;
            end else begin
              if (_T_88) begin
                out_valid_R_0 <= 1'h0;
              end
            end
          end else begin
            out_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_88) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      base_addr_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        if (_T_119) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            base_addr_R_taskID <= 10'h0;
          end else begin
            if (_T_119) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_119) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_119) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_119) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_119) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_119) begin
          base_addr_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            if (_T_119) begin
              base_addr_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_119) begin
            base_addr_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_126) begin
        if (_T_122) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_122) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_122) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_126) begin
        if (_T_122) begin
          idx_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            if (_T_122) begin
              idx_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_122) begin
            idx_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_126) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_127) begin
              state <= 1'h1;
            end
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_132) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UnTypLoad_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [9:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [9:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_165; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_168; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_5;
  reg [9:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_8;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_10;
  wire  _T_196; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_6; // @[LoadSimple.scala 81:27]
  wire [9:0] _GEN_7; // @[LoadSimple.scala 81:27]
  wire  _GEN_8; // @[LoadSimple.scala 81:27]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  _T_199; // @[HandShaking.scala 656:24]
  wire  _T_201; // @[HandShaking.scala 656:24]
  wire  _T_202; // @[HandShaking.scala 656:50]
  wire  _T_204; // @[HandShaking.scala 656:50]
  wire  complete; // @[HandShaking.scala 656:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_211; // @[Conditional.scala 37:30]
  wire  _T_212; // @[LoadSimple.scala 119:27]
  wire  _T_213; // @[LoadSimple.scala 120:31]
  wire [1:0] _GEN_10; // @[LoadSimple.scala 122:33]
  wire [1:0] _GEN_12; // @[LoadSimple.scala 120:45]
  wire  _GEN_14; // @[LoadSimple.scala 120:45]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire [1:0] _GEN_16; // @[LoadSimple.scala 119:44]
  wire  _GEN_18; // @[LoadSimple.scala 119:44]
  wire  _T_224; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_19; // @[LoadSimple.scala 135:30]
  wire  _GEN_21; // @[LoadSimple.scala 135:30]
  wire [1:0] _GEN_22; // @[LoadSimple.scala 135:30]
  wire  _T_234; // @[Conditional.scala 37:30]
  wire  _GEN_23; // @[LoadSimple.scala 149:22]
  wire  _GEN_25; // @[LoadSimple.scala 149:22]
  wire  _GEN_26; // @[LoadSimple.scala 149:22]
  wire [1:0] _GEN_27; // @[LoadSimple.scala 149:22]
  wire  _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  assign _T_165 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_165 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_165 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_168 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_168 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_168 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_168 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_196 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_196 ? io_GepAddr_bits_data : addr_R_data; // @[LoadSimple.scala 81:27]
  assign _GEN_7 = _T_196 ? io_GepAddr_bits_taskID : addr_R_taskID; // @[LoadSimple.scala 81:27]
  assign _GEN_8 = _T_196 ? io_GepAddr_bits_predicate : addr_R_predicate; // @[LoadSimple.scala 81:27]
  assign _GEN_9 = _T_196 ? 1'h1 : addr_valid_R; // @[LoadSimple.scala 81:27]
  assign _T_199 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_201 = _T_199 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_202 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_204 = _T_202 == 1'h0; // @[HandShaking.scala 656:50]
  assign complete = _T_201 | _T_204; // @[HandShaking.scala 656:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_211 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_212 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_213 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _GEN_10 = io_memReq_ready ? 2'h1 : state; // @[LoadSimple.scala 122:33]
  assign _GEN_12 = _T_213 ? _GEN_10 : 2'h2; // @[LoadSimple.scala 120:45]
  assign _GEN_14 = _T_213 ? _GEN_1 : 1'h1; // @[LoadSimple.scala 120:45]
  assign _GEN_15 = _T_212 ? _T_213 : 1'h0; // @[LoadSimple.scala 119:44]
  assign _GEN_16 = _T_212 ? _GEN_12 : state; // @[LoadSimple.scala 119:44]
  assign _GEN_18 = _T_212 ? _GEN_14 : _GEN_1; // @[LoadSimple.scala 119:44]
  assign _T_224 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _GEN_19 = io_memResp_valid ? io_memResp_data : data_R_data; // @[LoadSimple.scala 135:30]
  assign _GEN_21 = io_memResp_valid ? 1'h1 : _GEN_1; // @[LoadSimple.scala 135:30]
  assign _GEN_22 = io_memResp_valid ? 2'h2 : state; // @[LoadSimple.scala 135:30]
  assign _T_234 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_23 = complete ? 1'h0 : _GEN_9; // @[LoadSimple.scala 149:22]
  assign _GEN_25 = complete ? 1'h0 : _GEN_0; // @[LoadSimple.scala 149:22]
  assign _GEN_26 = complete ? 1'h0 : _GEN_2; // @[LoadSimple.scala 149:22]
  assign _GEN_27 = complete ? 2'h0 : state; // @[LoadSimple.scala 149:22]
  assign _GEN_28 = _T_234 ? _GEN_23 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_234 ? _GEN_25 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_234 ? _GEN_26 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_234 ? _GEN_27 : state; // @[Conditional.scala 39:67]
  assign _GEN_33 = _T_224 ? _GEN_19 : data_R_data; // @[Conditional.scala 39:67]
  assign _GEN_35 = _T_224 ? _GEN_21 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_224 ? _GEN_22 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_224 ? _GEN_9 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_224 ? _GEN_0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_40 = _T_224 ? _GEN_2 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_211 ? _GEN_16 : _GEN_36; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_211 ? _GEN_18 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_211 ? data_R_data : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_211 ? _GEN_9 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_211 ? _GEN_0 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_211 ? _GEN_2 : _GEN_40; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = addr_R_taskID | enable_R_taskID; // @[LoadSimple.scala 97:20 LoadSimple.scala 99:27]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_211 ? _GEN_15 : 1'h0; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_predicate = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_168) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_168) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_168) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_224) begin
          if (_T_168) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_168) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_168) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_165) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_224) begin
          if (_T_165) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_165) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_165) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_212) begin
          if (_T_213) begin
            if (_T_165) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_165) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_165) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_165) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_196) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 10'h0;
    end else begin
      if (_T_196) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_196) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_196) begin
          addr_valid_R <= 1'h1;
        end
      end else begin
        if (_T_224) begin
          if (_T_196) begin
            addr_valid_R <= 1'h1;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              if (_T_196) begin
                addr_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_196) begin
              addr_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_211)) begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_211) begin
        if (_T_212) begin
          if (_T_213) begin
            if (io_memReq_ready) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module FPMultiplier(
  input         clock,
  input  [31:0] io_dataa,
  input  [31:0] io_datab,
  output [31:0] io_result
);
  wire [31:0] fpmultiplier_result; // @[FPComputeNode.scala 245:28]
  wire [31:0] fpmultiplier_datab; // @[FPComputeNode.scala 245:28]
  wire [31:0] fpmultiplier_dataa; // @[FPComputeNode.scala 245:28]
  wire  fpmultiplier_clock; // @[FPComputeNode.scala 245:28]
  wire  fpmultiplier_clk_en; // @[FPComputeNode.scala 245:28]
  altfp_multiplier_11 fpmultiplier ( // @[FPComputeNode.scala 245:28]
    .result(fpmultiplier_result),
    .datab(fpmultiplier_datab),
    .dataa(fpmultiplier_dataa),
    .clock(fpmultiplier_clock),
    .clk_en(fpmultiplier_clk_en)
  );
  assign io_result = fpmultiplier_result; // @[FPComputeNode.scala 251:13]
  assign fpmultiplier_datab = io_datab; // @[FPComputeNode.scala 250:25]
  assign fpmultiplier_dataa = io_dataa; // @[FPComputeNode.scala 249:25]
  assign fpmultiplier_clock = clock; // @[FPComputeNode.scala 247:25]
  assign fpmultiplier_clk_en = 1'h1; // @[FPComputeNode.scala 248:26]
endmodule
module FPCustomMultiplierNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID,
  input  [31:0] io_RightIO_bits_data
);
  wire  FU_clock; // @[FPComputeNode.scala 551:18]
  wire [31:0] FU_io_dataa; // @[FPComputeNode.scala 551:18]
  wire [31:0] FU_io_datab; // @[FPComputeNode.scala 551:18]
  wire [31:0] FU_io_result; // @[FPComputeNode.scala 551:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[FPComputeNode.scala 527:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[FPComputeNode.scala 527:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[FPComputeNode.scala 528:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[FPComputeNode.scala 531:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[FPComputeNode.scala 531:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[FPComputeNode.scala 532:30]
  reg [31:0] _RAND_10;
  reg [9:0] out_data_R_taskID; // @[FPComputeNode.scala 537:27]
  reg [31:0] _RAND_11;
  reg [31:0] out_data_R_data; // @[FPComputeNode.scala 537:27]
  reg [31:0] _RAND_12;
  reg  state; // @[FPComputeNode.scala 540:22]
  reg [31:0] _RAND_13;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[FPComputeNode.scala 557:26]
  wire [31:0] _GEN_8; // @[FPComputeNode.scala 557:26]
  wire  _GEN_9; // @[FPComputeNode.scala 557:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[FPComputeNode.scala 563:27]
  wire [31:0] _GEN_12; // @[FPComputeNode.scala 563:27]
  wire  _GEN_13; // @[FPComputeNode.scala 563:27]
  wire  _T_119; // @[Conditional.scala 37:30]
  wire  _T_120; // @[FPComputeNode.scala 587:27]
  wire [9:0] _T_122; // @[FPComputeNode.scala 592:48]
  wire [9:0] _T_123; // @[FPComputeNode.scala 592:65]
  wire [31:0] _GEN_14; // @[FPComputeNode.scala 589:34]
  wire [9:0] _GEN_16; // @[FPComputeNode.scala 589:34]
  wire  _GEN_17; // @[FPComputeNode.scala 587:45]
  wire [31:0] _GEN_18; // @[FPComputeNode.scala 587:45]
  wire [9:0] _GEN_20; // @[FPComputeNode.scala 587:45]
  wire  _GEN_21; // @[FPComputeNode.scala 587:45]
  wire  _GEN_22; // @[FPComputeNode.scala 586:28]
  wire [31:0] _GEN_23; // @[FPComputeNode.scala 586:28]
  wire [9:0] _GEN_25; // @[FPComputeNode.scala 586:28]
  wire  _GEN_26; // @[FPComputeNode.scala 586:28]
  wire  _T_126; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[FPComputeNode.scala 599:26]
  wire  _GEN_28; // @[FPComputeNode.scala 599:26]
  wire  _GEN_29; // @[FPComputeNode.scala 599:26]
  wire  _GEN_31; // @[FPComputeNode.scala 599:26]
  wire  _GEN_32; // @[FPComputeNode.scala 599:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_40; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  FPMultiplier FU ( // @[FPComputeNode.scala 551:18]
    .clock(FU_clock),
    .io_dataa(FU_io_dataa),
    .io_datab(FU_io_datab),
    .io_result(FU_io_result)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[FPComputeNode.scala 557:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[FPComputeNode.scala 557:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[FPComputeNode.scala 557:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[FPComputeNode.scala 563:27]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[FPComputeNode.scala 563:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[FPComputeNode.scala 563:27]
  assign _T_119 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_120 = left_valid_R & right_valid_R; // @[FPComputeNode.scala 587:27]
  assign _T_122 = left_R_taskID | right_R_taskID; // @[FPComputeNode.scala 592:48]
  assign _T_123 = _T_122 | enable_R_taskID; // @[FPComputeNode.scala 592:65]
  assign _GEN_14 = enable_R_control ? FU_io_result : out_data_R_data; // @[FPComputeNode.scala 589:34]
  assign _GEN_16 = enable_R_control ? _T_123 : out_data_R_taskID; // @[FPComputeNode.scala 589:34]
  assign _GEN_17 = _T_120 ? 1'h1 : _GEN_1; // @[FPComputeNode.scala 587:45]
  assign _GEN_18 = _T_120 ? _GEN_14 : out_data_R_data; // @[FPComputeNode.scala 587:45]
  assign _GEN_20 = _T_120 ? _GEN_16 : out_data_R_taskID; // @[FPComputeNode.scala 587:45]
  assign _GEN_21 = _T_120 ? 1'h1 : state; // @[FPComputeNode.scala 587:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[FPComputeNode.scala 586:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : out_data_R_data; // @[FPComputeNode.scala 586:28]
  assign _GEN_25 = enable_valid_R ? _GEN_20 : out_data_R_taskID; // @[FPComputeNode.scala 586:28]
  assign _GEN_26 = enable_valid_R ? _GEN_21 : state; // @[FPComputeNode.scala 586:28]
  assign _T_126 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_126 ? 1'h0 : _GEN_9; // @[FPComputeNode.scala 599:26]
  assign _GEN_28 = _T_126 ? 1'h0 : _GEN_13; // @[FPComputeNode.scala 599:26]
  assign _GEN_29 = _T_126 ? 1'h0 : state; // @[FPComputeNode.scala 599:26]
  assign _GEN_31 = _T_126 ? 1'h0 : _GEN_0; // @[FPComputeNode.scala 599:26]
  assign _GEN_32 = _T_126 ? 1'h0 : _GEN_2; // @[FPComputeNode.scala 599:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_119 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_119 ? _GEN_23 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_42 = _T_119 ? _GEN_25 : out_data_R_taskID; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_119 ? _GEN_26 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_119 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_119 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_119 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_119 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = out_data_R_taskID; // @[FPComputeNode.scala 578:20]
  assign io_Out_0_bits_data = out_data_R_data; // @[FPComputeNode.scala 578:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[FPComputeNode.scala 556:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[FPComputeNode.scala 562:20]
  assign FU_clock = clock;
  assign FU_io_dataa = left_R_data; // @[FPComputeNode.scala 553:15]
  assign FU_io_datab = right_R_data; // @[FPComputeNode.scala 554:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_taskID = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_data_R_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_taskID <= 10'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            if (enable_R_control) begin
              out_data_R_taskID <= _T_123;
            end
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_result;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_3;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_4;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_5;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_6;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_7;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_8;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_9;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_8; // @[ComputeNode.scala 77:26]
  wire  _GEN_9; // @[ComputeNode.scala 77:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_12; // @[ComputeNode.scala 83:27]
  wire  _GEN_13; // @[ComputeNode.scala 83:27]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 110:34]
  wire  _GEN_17; // @[ComputeNode.scala 107:45]
  wire  _GEN_18; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_22; // @[ComputeNode.scala 106:28]
  wire  _GEN_23; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_24; // @[ComputeNode.scala 106:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[ComputeNode.scala 123:26]
  wire  _GEN_28; // @[ComputeNode.scala 123:26]
  wire  _GEN_29; // @[ComputeNode.scala 123:26]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[ComputeNode.scala 123:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[ComputeNode.scala 123:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  left_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  right_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  right_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_data_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module GepNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [9:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_1;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_2;
  reg  out_ready_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_1; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_5;
  wire  _T_98; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_100; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 186:29]
  wire  _GEN_3; // @[HandShaking.scala 186:29]
  wire  _T_103; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  wire  _GEN_6; // @[HandShaking.scala 197:27]
  reg [9:0] base_addr_R_taskID; // @[GepNode.scala 892:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 892:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 893:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 896:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 897:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 901:22]
  reg [31:0] _RAND_11;
  wire  _T_131; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_9; // @[GepNode.scala 917:31]
  wire [31:0] _GEN_10; // @[GepNode.scala 917:31]
  wire  _GEN_11; // @[GepNode.scala 917:31]
  wire  _T_134; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_14; // @[GepNode.scala 924:28]
  wire  _GEN_15; // @[GepNode.scala 924:28]
  wire [35:0] seek_value; // @[GepNode.scala 932:21]
  wire [35:0] _GEN_63; // @[GepNode.scala 940:35]
  wire [36:0] _T_137; // @[GepNode.scala 940:35]
  wire [35:0] data_out; // @[GepNode.scala 940:35]
  wire  _T_138; // @[Conditional.scala 37:30]
  wire  _T_139; // @[GepNode.scala 958:42]
  wire  _GEN_16; // @[GepNode.scala 958:64]
  wire  _GEN_17; // @[GepNode.scala 958:64]
  wire  _GEN_18; // @[GepNode.scala 958:64]
  wire  _GEN_19; // @[GepNode.scala 957:32]
  wire  _GEN_20; // @[GepNode.scala 957:32]
  wire  _GEN_21; // @[GepNode.scala 957:32]
  wire  _GEN_22; // @[GepNode.scala 956:28]
  wire  _GEN_23; // @[GepNode.scala 956:28]
  wire  _GEN_24; // @[GepNode.scala 956:28]
  wire  _T_147; // @[HandShaking.scala 222:83]
  wire  _T_148; // @[HandShaking.scala 222:83]
  wire  _T_149; // @[HandShaking.scala 224:11]
  wire [31:0] _GEN_25; // @[GepNode.scala 970:26]
  wire [31:0] _GEN_28; // @[GepNode.scala 970:26]
  wire [9:0] _GEN_29; // @[GepNode.scala 970:26]
  wire  _GEN_31; // @[GepNode.scala 970:26]
  wire  _GEN_32; // @[GepNode.scala 970:26]
  wire  _GEN_33; // @[GepNode.scala 970:26]
  wire  _GEN_34; // @[GepNode.scala 970:26]
  wire  _GEN_35; // @[GepNode.scala 970:26]
  wire  _GEN_36; // @[GepNode.scala 970:26]
  wire [31:0] _GEN_37; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_40; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_46; // @[Conditional.scala 39:67]
  wire  _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_48; // @[Conditional.scala 39:67]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  wire  _GEN_50; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_52; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_55; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_56; // @[Conditional.scala 40:58]
  wire  _GEN_58; // @[Conditional.scala 40:58]
  wire  _GEN_59; // @[Conditional.scala 40:58]
  wire  _GEN_60; // @[Conditional.scala 40:58]
  wire  _GEN_61; // @[Conditional.scala 40:58]
  wire  _GEN_62; // @[Conditional.scala 40:58]
  assign _T_98 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_98 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_98 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_100 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_100 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 186:29]
  assign _GEN_3 = _T_100 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 186:29]
  assign _T_103 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_103 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_6 = _T_103 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_131 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_131 ? io_baseAddress_bits_taskID : base_addr_R_taskID; // @[GepNode.scala 917:31]
  assign _GEN_10 = _T_131 ? io_baseAddress_bits_data : base_addr_R_data; // @[GepNode.scala 917:31]
  assign _GEN_11 = _T_131 ? 1'h1 : base_addr_valid_R; // @[GepNode.scala 917:31]
  assign _T_134 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_14 = _T_134 ? io_idx_0_bits_data : idx_R_0_data; // @[GepNode.scala 924:28]
  assign _GEN_15 = _T_134 ? 1'h1 : idx_valid_R_0; // @[GepNode.scala 924:28]
  assign seek_value = idx_R_0_data * 32'h8; // @[GepNode.scala 932:21]
  assign _GEN_63 = {{4'd0}, base_addr_R_data}; // @[GepNode.scala 940:35]
  assign _T_137 = _GEN_63 + seek_value; // @[GepNode.scala 940:35]
  assign data_out = _GEN_63 + seek_value; // @[GepNode.scala 940:35]
  assign _T_138 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_139 = idx_valid_R_0 & base_addr_valid_R; // @[GepNode.scala 958:42]
  assign _GEN_16 = _T_139 ? 1'h1 : _GEN_1; // @[GepNode.scala 958:64]
  assign _GEN_17 = _T_139 ? 1'h1 : _GEN_3; // @[GepNode.scala 958:64]
  assign _GEN_18 = _T_139 ? 1'h1 : state; // @[GepNode.scala 958:64]
  assign _GEN_19 = enable_R_control ? _GEN_16 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_20 = enable_R_control ? _GEN_17 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_21 = enable_R_control ? _GEN_18 : 1'h1; // @[GepNode.scala 957:32]
  assign _GEN_22 = enable_valid_R ? _GEN_19 : _GEN_1; // @[GepNode.scala 956:28]
  assign _GEN_23 = enable_valid_R ? _GEN_20 : _GEN_3; // @[GepNode.scala 956:28]
  assign _GEN_24 = enable_valid_R ? _GEN_21 : state; // @[GepNode.scala 956:28]
  assign _T_147 = out_ready_R_0 | _T_98; // @[HandShaking.scala 222:83]
  assign _T_148 = out_ready_R_1 | _T_100; // @[HandShaking.scala 222:83]
  assign _T_149 = _T_147 & _T_148; // @[HandShaking.scala 224:11]
  assign _GEN_25 = _T_149 ? 32'h0 : _GEN_14; // @[GepNode.scala 970:26]
  assign _GEN_28 = _T_149 ? 32'h0 : _GEN_10; // @[GepNode.scala 970:26]
  assign _GEN_29 = _T_149 ? 10'h0 : _GEN_9; // @[GepNode.scala 970:26]
  assign _GEN_31 = _T_149 ? 1'h0 : _GEN_15; // @[GepNode.scala 970:26]
  assign _GEN_32 = _T_149 ? 1'h0 : _GEN_11; // @[GepNode.scala 970:26]
  assign _GEN_33 = _T_149 ? 1'h0 : state; // @[GepNode.scala 970:26]
  assign _GEN_34 = _T_149 ? 1'h0 : _GEN_0; // @[GepNode.scala 970:26]
  assign _GEN_35 = _T_149 ? 1'h0 : _GEN_2; // @[GepNode.scala 970:26]
  assign _GEN_36 = _T_149 ? 1'h0 : _GEN_4; // @[GepNode.scala 970:26]
  assign _GEN_37 = state ? _GEN_25 : _GEN_14; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_28 : _GEN_10; // @[Conditional.scala 39:67]
  assign _GEN_41 = state ? _GEN_29 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_31 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_44 = state ? _GEN_32 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_45 = state ? _GEN_33 : state; // @[Conditional.scala 39:67]
  assign _GEN_46 = state ? _GEN_34 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_47 = state ? _GEN_35 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_48 = state ? _GEN_36 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_49 = _T_138 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_138 ? _GEN_23 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_138 ? _GEN_24 : _GEN_45; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_138 ? _GEN_14 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_138 ? _GEN_10 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_56 = _T_138 ? _GEN_9 : _GEN_41; // @[Conditional.scala 40:58]
  assign _GEN_58 = _T_138 ? _GEN_15 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_59 = _T_138 ? _GEN_11 : _GEN_44; // @[Conditional.scala 40:58]
  assign _GEN_60 = _T_138 ? _GEN_0 : _GEN_46; // @[Conditional.scala 40:58]
  assign _GEN_61 = _T_138 ? _GEN_2 : _GEN_47; // @[Conditional.scala 40:58]
  assign _GEN_62 = _T_138 ? _GEN_4 : _GEN_48; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 945:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 946:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 944:25]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 184:21]
  assign io_Out_1_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 946:27]
  assign io_Out_1_bits_data = data_out[31:0]; // @[GepNode.scala 944:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 916:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 923:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_control = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_103) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_138) begin
        if (_T_103) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_103) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_103) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_138) begin
        if (_T_98) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_98) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_98) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_138) begin
        if (_T_100) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_100) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_100) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_138) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_139) begin
              out_valid_R_0 <= 1'h1;
            end else begin
              if (_T_98) begin
                out_valid_R_0 <= 1'h0;
              end
            end
          end else begin
            out_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_98) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_98) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_138) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_139) begin
              out_valid_R_1 <= 1'h1;
            end else begin
              if (_T_100) begin
                out_valid_R_1 <= 1'h0;
              end
            end
          end else begin
            out_valid_R_1 <= 1'h1;
          end
        end else begin
          if (_T_100) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_100) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      base_addr_R_taskID <= 10'h0;
    end else begin
      if (_T_138) begin
        if (_T_131) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            base_addr_R_taskID <= 10'h0;
          end else begin
            if (_T_131) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_131) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_138) begin
        if (_T_131) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_131) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_131) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_138) begin
        if (_T_131) begin
          base_addr_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            if (_T_131) begin
              base_addr_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_131) begin
            base_addr_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_138) begin
        if (_T_134) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_134) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_134) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_138) begin
        if (_T_134) begin
          idx_valid_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            if (_T_134) begin
              idx_valid_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_134) begin
            idx_valid_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_138) begin
        if (enable_valid_R) begin
          if (enable_R_control) begin
            if (_T_139) begin
              state <= 1'h1;
            end
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UnTypLoad_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [9:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [9:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 538:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 539:28]
  reg [31:0] _RAND_4;
  wire  _T_165; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 565:29]
  wire  _GEN_1; // @[HandShaking.scala 565:29]
  wire  _T_168; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_5;
  reg [9:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_8;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_10;
  wire  _T_196; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_6; // @[LoadSimple.scala 81:27]
  wire [9:0] _GEN_7; // @[LoadSimple.scala 81:27]
  wire  _GEN_8; // @[LoadSimple.scala 81:27]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  _T_199; // @[HandShaking.scala 656:24]
  wire  _T_201; // @[HandShaking.scala 656:24]
  wire  _T_202; // @[HandShaking.scala 656:50]
  wire  _T_204; // @[HandShaking.scala 656:50]
  wire  complete; // @[HandShaking.scala 656:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_211; // @[Conditional.scala 37:30]
  wire  _T_212; // @[LoadSimple.scala 119:27]
  wire  _T_213; // @[LoadSimple.scala 120:31]
  wire [1:0] _GEN_10; // @[LoadSimple.scala 122:33]
  wire [1:0] _GEN_12; // @[LoadSimple.scala 120:45]
  wire  _GEN_14; // @[LoadSimple.scala 120:45]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire [1:0] _GEN_16; // @[LoadSimple.scala 119:44]
  wire  _GEN_18; // @[LoadSimple.scala 119:44]
  wire  _T_224; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_19; // @[LoadSimple.scala 135:30]
  wire  _GEN_21; // @[LoadSimple.scala 135:30]
  wire [1:0] _GEN_22; // @[LoadSimple.scala 135:30]
  wire  _T_234; // @[Conditional.scala 37:30]
  wire  _GEN_23; // @[LoadSimple.scala 149:22]
  wire  _GEN_25; // @[LoadSimple.scala 149:22]
  wire  _GEN_26; // @[LoadSimple.scala 149:22]
  wire [1:0] _GEN_27; // @[LoadSimple.scala 149:22]
  wire  _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  assign _T_165 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_165 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 565:29]
  assign _GEN_1 = _T_165 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 565:29]
  assign _T_168 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_168 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_168 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_168 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_196 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_196 ? io_GepAddr_bits_data : addr_R_data; // @[LoadSimple.scala 81:27]
  assign _GEN_7 = _T_196 ? io_GepAddr_bits_taskID : addr_R_taskID; // @[LoadSimple.scala 81:27]
  assign _GEN_8 = _T_196 ? io_GepAddr_bits_predicate : addr_R_predicate; // @[LoadSimple.scala 81:27]
  assign _GEN_9 = _T_196 ? 1'h1 : addr_valid_R; // @[LoadSimple.scala 81:27]
  assign _T_199 = ~ out_ready_R_0; // @[HandShaking.scala 656:24]
  assign _T_201 = _T_199 == 1'h0; // @[HandShaking.scala 656:24]
  assign _T_202 = ~ io_Out_0_ready; // @[HandShaking.scala 656:50]
  assign _T_204 = _T_202 == 1'h0; // @[HandShaking.scala 656:50]
  assign complete = _T_201 | _T_204; // @[HandShaking.scala 656:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_211 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_212 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_213 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _GEN_10 = io_memReq_ready ? 2'h1 : state; // @[LoadSimple.scala 122:33]
  assign _GEN_12 = _T_213 ? _GEN_10 : 2'h2; // @[LoadSimple.scala 120:45]
  assign _GEN_14 = _T_213 ? _GEN_1 : 1'h1; // @[LoadSimple.scala 120:45]
  assign _GEN_15 = _T_212 ? _T_213 : 1'h0; // @[LoadSimple.scala 119:44]
  assign _GEN_16 = _T_212 ? _GEN_12 : state; // @[LoadSimple.scala 119:44]
  assign _GEN_18 = _T_212 ? _GEN_14 : _GEN_1; // @[LoadSimple.scala 119:44]
  assign _T_224 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _GEN_19 = io_memResp_valid ? io_memResp_data : data_R_data; // @[LoadSimple.scala 135:30]
  assign _GEN_21 = io_memResp_valid ? 1'h1 : _GEN_1; // @[LoadSimple.scala 135:30]
  assign _GEN_22 = io_memResp_valid ? 2'h2 : state; // @[LoadSimple.scala 135:30]
  assign _T_234 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_23 = complete ? 1'h0 : _GEN_9; // @[LoadSimple.scala 149:22]
  assign _GEN_25 = complete ? 1'h0 : _GEN_0; // @[LoadSimple.scala 149:22]
  assign _GEN_26 = complete ? 1'h0 : _GEN_2; // @[LoadSimple.scala 149:22]
  assign _GEN_27 = complete ? 2'h0 : state; // @[LoadSimple.scala 149:22]
  assign _GEN_28 = _T_234 ? _GEN_23 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_234 ? _GEN_25 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_234 ? _GEN_26 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_234 ? _GEN_27 : state; // @[Conditional.scala 39:67]
  assign _GEN_33 = _T_224 ? _GEN_19 : data_R_data; // @[Conditional.scala 39:67]
  assign _GEN_35 = _T_224 ? _GEN_21 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_224 ? _GEN_22 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_37 = _T_224 ? _GEN_9 : _GEN_28; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_224 ? _GEN_0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_40 = _T_224 ? _GEN_2 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_211 ? _GEN_16 : _GEN_36; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_211 ? _GEN_18 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_211 ? data_R_data : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_211 ? _GEN_9 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_211 ? _GEN_0 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_211 ? _GEN_2 : _GEN_40; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 563:21]
  assign io_Out_0_bits_taskID = addr_R_taskID | enable_R_taskID; // @[LoadSimple.scala 97:20 LoadSimple.scala 99:27]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_211 ? _GEN_15 : 1'h0; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_predicate = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_168) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_168) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_168) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_224) begin
          if (_T_168) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_168) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_168) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_165) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_224) begin
          if (_T_165) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_165) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_165) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_212) begin
          if (_T_213) begin
            if (_T_165) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_165) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_165) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_165) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_196) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 10'h0;
    end else begin
      if (_T_196) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_196) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_211) begin
        if (_T_196) begin
          addr_valid_R <= 1'h1;
        end
      end else begin
        if (_T_224) begin
          if (_T_196) begin
            addr_valid_R <= 1'h1;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              if (_T_196) begin
                addr_valid_R <= 1'h1;
              end
            end
          end else begin
            if (_T_196) begin
              addr_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_211)) begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_211) begin
        if (_T_212) begin
          if (_T_213) begin
            if (io_memReq_ready) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_224) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_234) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module FPAdder(
  input         clock,
  input  [31:0] io_dataa,
  input  [31:0] io_datab,
  output [31:0] io_result
);
  wire [31:0] fpadder_result; // @[FPComputeNode.scala 211:23]
  wire [31:0] fpadder_datab; // @[FPComputeNode.scala 211:23]
  wire [31:0] fpadder_dataa; // @[FPComputeNode.scala 211:23]
  wire  fpadder_clock; // @[FPComputeNode.scala 211:23]
  wire  fpadder_clk_en; // @[FPComputeNode.scala 211:23]
  altfp_adder_13 fpadder ( // @[FPComputeNode.scala 211:23]
    .result(fpadder_result),
    .datab(fpadder_datab),
    .dataa(fpadder_dataa),
    .clock(fpadder_clock),
    .clk_en(fpadder_clk_en)
  );
  assign io_result = fpadder_result; // @[FPComputeNode.scala 217:13]
  assign fpadder_datab = io_datab; // @[FPComputeNode.scala 216:20]
  assign fpadder_dataa = io_dataa; // @[FPComputeNode.scala 215:20]
  assign fpadder_clock = clock; // @[FPComputeNode.scala 213:20]
  assign fpadder_clk_en = 1'h1; // @[FPComputeNode.scala 214:21]
endmodule
module FPCustomAdderNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID,
  input  [31:0] io_RightIO_bits_data
);
  wire  FU_clock; // @[FPComputeNode.scala 320:18]
  wire [31:0] FU_io_dataa; // @[FPComputeNode.scala 320:18]
  wire [31:0] FU_io_datab; // @[FPComputeNode.scala 320:18]
  wire [31:0] FU_io_result; // @[FPComputeNode.scala 320:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[FPComputeNode.scala 296:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[FPComputeNode.scala 296:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[FPComputeNode.scala 297:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[FPComputeNode.scala 300:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[FPComputeNode.scala 300:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[FPComputeNode.scala 301:30]
  reg [31:0] _RAND_10;
  reg [9:0] out_data_R_taskID; // @[FPComputeNode.scala 306:27]
  reg [31:0] _RAND_11;
  reg [31:0] out_data_R_data; // @[FPComputeNode.scala 306:27]
  reg [31:0] _RAND_12;
  reg  state; // @[FPComputeNode.scala 309:22]
  reg [31:0] _RAND_13;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[FPComputeNode.scala 326:26]
  wire [31:0] _GEN_8; // @[FPComputeNode.scala 326:26]
  wire  _GEN_9; // @[FPComputeNode.scala 326:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[FPComputeNode.scala 332:27]
  wire [31:0] _GEN_12; // @[FPComputeNode.scala 332:27]
  wire  _GEN_13; // @[FPComputeNode.scala 332:27]
  wire  _T_119; // @[Conditional.scala 37:30]
  wire  _T_120; // @[FPComputeNode.scala 356:27]
  wire [9:0] _T_122; // @[FPComputeNode.scala 361:48]
  wire [9:0] _T_123; // @[FPComputeNode.scala 361:65]
  wire [31:0] _GEN_14; // @[FPComputeNode.scala 358:34]
  wire [9:0] _GEN_16; // @[FPComputeNode.scala 358:34]
  wire  _GEN_17; // @[FPComputeNode.scala 356:45]
  wire [31:0] _GEN_18; // @[FPComputeNode.scala 356:45]
  wire [9:0] _GEN_20; // @[FPComputeNode.scala 356:45]
  wire  _GEN_21; // @[FPComputeNode.scala 356:45]
  wire  _GEN_22; // @[FPComputeNode.scala 355:28]
  wire [31:0] _GEN_23; // @[FPComputeNode.scala 355:28]
  wire [9:0] _GEN_25; // @[FPComputeNode.scala 355:28]
  wire  _GEN_26; // @[FPComputeNode.scala 355:28]
  wire  _T_126; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[FPComputeNode.scala 368:26]
  wire  _GEN_28; // @[FPComputeNode.scala 368:26]
  wire  _GEN_29; // @[FPComputeNode.scala 368:26]
  wire  _GEN_31; // @[FPComputeNode.scala 368:26]
  wire  _GEN_32; // @[FPComputeNode.scala 368:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_40; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_42; // @[Conditional.scala 40:58]
  wire  _GEN_43; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  FPAdder FU ( // @[FPComputeNode.scala 320:18]
    .clock(FU_clock),
    .io_dataa(FU_io_dataa),
    .io_datab(FU_io_datab),
    .io_result(FU_io_result)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[FPComputeNode.scala 326:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[FPComputeNode.scala 326:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[FPComputeNode.scala 326:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[FPComputeNode.scala 332:27]
  assign _GEN_12 = _T_117 ? io_RightIO_bits_data : right_R_data; // @[FPComputeNode.scala 332:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[FPComputeNode.scala 332:27]
  assign _T_119 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_120 = left_valid_R & right_valid_R; // @[FPComputeNode.scala 356:27]
  assign _T_122 = left_R_taskID | right_R_taskID; // @[FPComputeNode.scala 361:48]
  assign _T_123 = _T_122 | enable_R_taskID; // @[FPComputeNode.scala 361:65]
  assign _GEN_14 = enable_R_control ? FU_io_result : out_data_R_data; // @[FPComputeNode.scala 358:34]
  assign _GEN_16 = enable_R_control ? _T_123 : out_data_R_taskID; // @[FPComputeNode.scala 358:34]
  assign _GEN_17 = _T_120 ? 1'h1 : _GEN_1; // @[FPComputeNode.scala 356:45]
  assign _GEN_18 = _T_120 ? _GEN_14 : out_data_R_data; // @[FPComputeNode.scala 356:45]
  assign _GEN_20 = _T_120 ? _GEN_16 : out_data_R_taskID; // @[FPComputeNode.scala 356:45]
  assign _GEN_21 = _T_120 ? 1'h1 : state; // @[FPComputeNode.scala 356:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[FPComputeNode.scala 355:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : out_data_R_data; // @[FPComputeNode.scala 355:28]
  assign _GEN_25 = enable_valid_R ? _GEN_20 : out_data_R_taskID; // @[FPComputeNode.scala 355:28]
  assign _GEN_26 = enable_valid_R ? _GEN_21 : state; // @[FPComputeNode.scala 355:28]
  assign _T_126 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_126 ? 1'h0 : _GEN_9; // @[FPComputeNode.scala 368:26]
  assign _GEN_28 = _T_126 ? 1'h0 : _GEN_13; // @[FPComputeNode.scala 368:26]
  assign _GEN_29 = _T_126 ? 1'h0 : state; // @[FPComputeNode.scala 368:26]
  assign _GEN_31 = _T_126 ? 1'h0 : _GEN_0; // @[FPComputeNode.scala 368:26]
  assign _GEN_32 = _T_126 ? 1'h0 : _GEN_2; // @[FPComputeNode.scala 368:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_119 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_119 ? _GEN_23 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_42 = _T_119 ? _GEN_25 : out_data_R_taskID; // @[Conditional.scala 40:58]
  assign _GEN_43 = _T_119 ? _GEN_26 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_119 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_119 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_119 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_119 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = out_data_R_taskID; // @[FPComputeNode.scala 347:20]
  assign io_Out_0_bits_data = out_data_R_data; // @[FPComputeNode.scala 347:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[FPComputeNode.scala 325:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[FPComputeNode.scala 331:20]
  assign FU_clock = clock;
  assign FU_io_dataa = left_R_data; // @[FPComputeNode.scala 322:15]
  assign FU_io_datab = right_R_data; // @[FPComputeNode.scala 323:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_taskID = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_data_R_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_119) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_taskID <= 10'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            if (enable_R_control) begin
              out_data_R_taskID <= _T_123;
            end
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_result;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_119) begin
        if (enable_valid_R) begin
          if (_T_120) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_126) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UnTypStore(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [9:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [9:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [9:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 525:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 526:31]
  reg [31:0] _RAND_2;
  wire  _T_180; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 584:27]
  wire  _GEN_3; // @[HandShaking.scala 584:27]
  wire [9:0] _GEN_4; // @[HandShaking.scala 584:27]
  reg [9:0] addr_R_taskID; // @[StoreSimple.scala 63:23]
  reg [31:0] _RAND_3;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 63:23]
  reg [31:0] _RAND_4;
  reg [9:0] data_R_taskID; // @[StoreSimple.scala 64:23]
  reg [31:0] _RAND_5;
  reg [31:0] data_R_data; // @[StoreSimple.scala 64:23]
  reg [31:0] _RAND_6;
  reg  addr_valid_R; // @[StoreSimple.scala 65:29]
  reg [31:0] _RAND_7;
  reg  data_valid_R; // @[StoreSimple.scala 66:29]
  reg [31:0] _RAND_8;
  reg [1:0] state; // @[StoreSimple.scala 70:22]
  reg [31:0] _RAND_9;
  wire  _T_212; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_6; // @[StoreSimple.scala 91:27]
  wire [9:0] _GEN_7; // @[StoreSimple.scala 91:27]
  wire  _GEN_9; // @[StoreSimple.scala 91:27]
  wire  _T_215; // @[Decoupled.scala 37:37]
  wire [31:0] _GEN_10; // @[StoreSimple.scala 99:26]
  wire [9:0] _GEN_11; // @[StoreSimple.scala 99:26]
  wire  _GEN_13; // @[StoreSimple.scala 99:26]
  wire [9:0] _T_217; // @[StoreSimple.scala 108:44]
  wire  mem_req_fire; // @[StoreSimple.scala 122:51]
  wire  _T_234; // @[Conditional.scala 37:30]
  wire  _T_235; // @[StoreSimple.scala 128:27]
  wire  _T_236; // @[StoreSimple.scala 129:33]
  wire [1:0] _GEN_14; // @[StoreSimple.scala 131:35]
  wire [1:0] _GEN_16; // @[StoreSimple.scala 129:50]
  wire  _GEN_19; // @[StoreSimple.scala 128:44]
  wire [1:0] _GEN_20; // @[StoreSimple.scala 128:44]
  wire  _GEN_23; // @[StoreSimple.scala 127:28]
  wire [1:0] _GEN_24; // @[StoreSimple.scala 127:28]
  wire  _T_247; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_28; // @[StoreSimple.scala 144:30]
  wire  _T_256; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_40; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_44; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_45; // @[Conditional.scala 39:67]
  wire  _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_49; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_50; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_52; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_53; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_56; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_57; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_60; // @[Conditional.scala 39:67]
  wire  _GEN_62; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_64; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_67; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_68; // @[Conditional.scala 40:58]
  wire  _GEN_70; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_71; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_72; // @[Conditional.scala 40:58]
  wire  _GEN_73; // @[Conditional.scala 40:58]
  wire  _GEN_75; // @[Conditional.scala 40:58]
  assign _T_180 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_180 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 584:27]
  assign _GEN_3 = _T_180 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 584:27]
  assign _GEN_4 = _T_180 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 584:27]
  assign _T_212 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_212 ? io_GepAddr_bits_data : addr_R_data; // @[StoreSimple.scala 91:27]
  assign _GEN_7 = _T_212 ? io_GepAddr_bits_taskID : addr_R_taskID; // @[StoreSimple.scala 91:27]
  assign _GEN_9 = _T_212 ? 1'h1 : addr_valid_R; // @[StoreSimple.scala 91:27]
  assign _T_215 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 37:37]
  assign _GEN_10 = _T_215 ? io_inData_bits_data : data_R_data; // @[StoreSimple.scala 99:26]
  assign _GEN_11 = _T_215 ? io_inData_bits_taskID : data_R_taskID; // @[StoreSimple.scala 99:26]
  assign _GEN_13 = _T_215 ? 1'h1 : data_valid_R; // @[StoreSimple.scala 99:26]
  assign _T_217 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 108:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 122:51]
  assign _T_234 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_235 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 128:27]
  assign _T_236 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 129:33]
  assign _GEN_14 = io_memReq_ready ? 2'h1 : state; // @[StoreSimple.scala 131:35]
  assign _GEN_16 = _T_236 ? _GEN_14 : 2'h2; // @[StoreSimple.scala 129:50]
  assign _GEN_19 = _T_235 ? _T_236 : 1'h0; // @[StoreSimple.scala 128:44]
  assign _GEN_20 = _T_235 ? _GEN_16 : state; // @[StoreSimple.scala 128:44]
  assign _GEN_23 = enable_valid_R ? _GEN_19 : 1'h0; // @[StoreSimple.scala 127:28]
  assign _GEN_24 = enable_valid_R ? _GEN_20 : state; // @[StoreSimple.scala 127:28]
  assign _T_247 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _GEN_28 = io_memResp_valid ? 2'h2 : state; // @[StoreSimple.scala 144:30]
  assign _T_256 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_40 = _T_256 ? 32'h0 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_256 ? 10'h0 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_256 ? 1'h0 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_44 = _T_256 ? 32'h0 : _GEN_10; // @[Conditional.scala 39:67]
  assign _GEN_45 = _T_256 ? 10'h0 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_47 = _T_256 ? 1'h0 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_49 = _T_256 ? 1'h0 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_50 = _T_256 ? 2'h0 : state; // @[Conditional.scala 39:67]
  assign _GEN_52 = _T_247 ? _GEN_28 : _GEN_50; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_247 ? _GEN_6 : _GEN_40; // @[Conditional.scala 39:67]
  assign _GEN_54 = _T_247 ? _GEN_7 : _GEN_41; // @[Conditional.scala 39:67]
  assign _GEN_56 = _T_247 ? _GEN_9 : _GEN_43; // @[Conditional.scala 39:67]
  assign _GEN_57 = _T_247 ? _GEN_10 : _GEN_44; // @[Conditional.scala 39:67]
  assign _GEN_58 = _T_247 ? _GEN_11 : _GEN_45; // @[Conditional.scala 39:67]
  assign _GEN_60 = _T_247 ? _GEN_13 : _GEN_47; // @[Conditional.scala 39:67]
  assign _GEN_62 = _T_247 ? _GEN_2 : _GEN_49; // @[Conditional.scala 39:67]
  assign _GEN_64 = _T_234 ? _GEN_24 : _GEN_52; // @[Conditional.scala 40:58]
  assign _GEN_67 = _T_234 ? _GEN_6 : _GEN_53; // @[Conditional.scala 40:58]
  assign _GEN_68 = _T_234 ? _GEN_7 : _GEN_54; // @[Conditional.scala 40:58]
  assign _GEN_70 = _T_234 ? _GEN_9 : _GEN_56; // @[Conditional.scala 40:58]
  assign _GEN_71 = _T_234 ? _GEN_10 : _GEN_57; // @[Conditional.scala 40:58]
  assign _GEN_72 = _T_234 ? _GEN_11 : _GEN_58; // @[Conditional.scala 40:58]
  assign _GEN_73 = _T_234 ? _GEN_13 : _GEN_60; // @[Conditional.scala 40:58]
  assign _GEN_75 = _T_234 ? _GEN_2 : _GEN_62; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 583:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 86:20 StoreSimple.scala 90:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 87:19]
  assign io_memReq_valid = _T_234 ? _GEN_23 : 1'h0; // @[StoreSimple.scala 117:19 StoreSimple.scala 130:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 111:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 112:23]
  assign io_memReq_bits_taskID = _T_217 | enable_R_taskID; // @[StoreSimple.scala 115:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  addr_R_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  data_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  data_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_180) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_180) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_234) begin
        if (_T_180) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_247) begin
          if (_T_180) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_256) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_180) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_taskID <= 10'h0;
    end else begin
      if (_T_234) begin
        if (_T_212) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_247) begin
          if (_T_212) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_256) begin
            addr_R_taskID <= 10'h0;
          end else begin
            if (_T_212) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_234) begin
        if (_T_212) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_247) begin
          if (_T_212) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_256) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_212) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 10'h0;
    end else begin
      if (_T_234) begin
        if (_T_215) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_247) begin
          if (_T_215) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_256) begin
            data_R_taskID <= 10'h0;
          end else begin
            if (_T_215) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_234) begin
        if (_T_215) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_247) begin
          if (_T_215) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_256) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_215) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_234) begin
        if (_T_212) begin
          addr_valid_R <= 1'h1;
        end
      end else begin
        if (_T_247) begin
          if (_T_212) begin
            addr_valid_R <= 1'h1;
          end
        end else begin
          if (_T_256) begin
            addr_valid_R <= 1'h0;
          end else begin
            if (_T_212) begin
              addr_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_234) begin
        if (_T_215) begin
          data_valid_R <= 1'h1;
        end
      end else begin
        if (_T_247) begin
          if (_T_215) begin
            data_valid_R <= 1'h1;
          end
        end else begin
          if (_T_256) begin
            data_valid_R <= 1'h0;
          end else begin
            if (_T_215) begin
              data_valid_R <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_234) begin
        if (enable_valid_R) begin
          if (_T_235) begin
            if (_T_236) begin
              if (io_memReq_ready) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_247) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_256) begin
            state <= 2'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_6;
  wire  _T_86; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 186:29]
  wire  _GEN_3; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_5; // @[HandShaking.scala 197:27]
  wire  _GEN_6; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_7;
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_9;
  reg [9:0] right_R_taskID; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_10;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_11;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_14;
  wire  _T_126; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_9; // @[ComputeNode.scala 77:26]
  wire [31:0] _GEN_10; // @[ComputeNode.scala 77:26]
  wire  _GEN_11; // @[ComputeNode.scala 77:26]
  wire  _T_129; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_13; // @[ComputeNode.scala 83:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 83:27]
  wire  _GEN_15; // @[ComputeNode.scala 83:27]
  wire [9:0] _T_131; // @[ComputeNode.scala 98:44]
  wire  _T_135; // @[Conditional.scala 37:30]
  wire  _T_136; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 110:34]
  wire  _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_20; // @[ComputeNode.scala 107:45]
  wire  _GEN_21; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_22; // @[ComputeNode.scala 107:45]
  wire  _GEN_25; // @[ComputeNode.scala 106:28]
  wire  _GEN_26; // @[ComputeNode.scala 106:28]
  wire  _GEN_27; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_28; // @[ComputeNode.scala 106:28]
  wire  _T_147; // @[HandShaking.scala 222:83]
  wire  _T_148; // @[HandShaking.scala 222:83]
  wire  _T_149; // @[HandShaking.scala 224:11]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[ComputeNode.scala 123:26]
  wire  _GEN_35; // @[ComputeNode.scala 123:26]
  wire  _GEN_36; // @[ComputeNode.scala 123:26]
  wire  _GEN_37; // @[ComputeNode.scala 123:26]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire  _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_86 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_86 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_86 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_88 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_88 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 186:29]
  assign _GEN_3 = _T_88 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_5 = _T_91 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_6 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_126 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_126 ? io_LeftIO_bits_taskID : left_R_taskID; // @[ComputeNode.scala 77:26]
  assign _GEN_10 = _T_126 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_11 = _T_126 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_129 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_13 = _T_129 ? io_RightIO_bits_taskID : right_R_taskID; // @[ComputeNode.scala 83:27]
  assign _GEN_14 = _T_129 ? 32'h1 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_15 = _T_129 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_131 = left_R_taskID | right_R_taskID; // @[ComputeNode.scala 98:44]
  assign _T_135 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_136 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_16 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_19 = _T_136 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_20 = _T_136 ? 1'h1 : _GEN_3; // @[ComputeNode.scala 107:45]
  assign _GEN_21 = _T_136 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = _T_136 ? _GEN_16 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_25 = enable_valid_R ? _GEN_19 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_26 = enable_valid_R ? _GEN_20 : _GEN_3; // @[ComputeNode.scala 106:28]
  assign _GEN_27 = enable_valid_R ? _GEN_21 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_28 = enable_valid_R ? _GEN_22 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_147 = out_ready_R_0 | _T_86; // @[HandShaking.scala 222:83]
  assign _T_148 = out_ready_R_1 | _T_88; // @[HandShaking.scala 222:83]
  assign _T_149 = _T_147 & _T_148; // @[HandShaking.scala 224:11]
  assign _GEN_31 = _T_149 ? 1'h0 : _GEN_11; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_149 ? 1'h0 : _GEN_15; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = _T_149 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_35 = _T_149 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_36 = _T_149 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_37 = _T_149 ? 1'h0 : _GEN_4; // @[ComputeNode.scala 123:26]
  assign _GEN_38 = state ? _GEN_31 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_32 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_33 : state; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_35 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_36 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_44 = state ? _GEN_37 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_45 = _T_135 ? _GEN_25 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_135 ? _GEN_26 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_135 ? _GEN_27 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_135 ? _GEN_28 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_135 ? _GEN_11 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_135 ? _GEN_15 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_135 ? _GEN_0 : _GEN_42; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_135 ? _GEN_2 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_135 ? _GEN_4 : _GEN_44; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 184:21]
  assign io_Out_1_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_1_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_R_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_valid_R = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_91) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_86) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_86) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_86) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_88) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_86) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_86) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_86) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_1 <= 1'h1;
          end else begin
            if (_T_88) begin
              out_valid_R_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_88) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_126) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_126) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_126) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_129) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_129) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_129) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_129) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_129) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UCMP(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire  _T_11; // @[Comparision.scala 81:32]
  assign _T_11 = io_in1 == io_in2; // @[Comparision.scala 81:32]
  assign io_out = {{31'd0}, _T_11}; // @[Comparision.scala 90:10]
endmodule
module IcmpNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_in2; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_out; // @[IcmpNode.scala 192:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[IcmpNode.scala 170:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[IcmpNode.scala 174:30]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R_data; // @[IcmpNode.scala 179:27]
  reg [31:0] _RAND_11;
  reg  state; // @[IcmpNode.scala 182:22]
  reg [31:0] _RAND_12;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[IcmpNode.scala 197:26]
  wire [31:0] _GEN_8; // @[IcmpNode.scala 197:26]
  wire  _GEN_9; // @[IcmpNode.scala 197:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[IcmpNode.scala 203:27]
  wire [31:0] _GEN_12; // @[IcmpNode.scala 203:27]
  wire  _GEN_13; // @[IcmpNode.scala 203:27]
  wire [9:0] _T_119; // @[IcmpNode.scala 218:44]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[IcmpNode.scala 227:27]
  wire [31:0] _GEN_14; // @[IcmpNode.scala 230:34]
  wire  _GEN_17; // @[IcmpNode.scala 227:45]
  wire  _GEN_18; // @[IcmpNode.scala 227:45]
  wire [31:0] _GEN_19; // @[IcmpNode.scala 227:45]
  wire  _GEN_22; // @[IcmpNode.scala 226:28]
  wire  _GEN_23; // @[IcmpNode.scala 226:28]
  wire [31:0] _GEN_24; // @[IcmpNode.scala 226:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[IcmpNode.scala 247:26]
  wire  _GEN_28; // @[IcmpNode.scala 247:26]
  wire  _GEN_29; // @[IcmpNode.scala 247:26]
  wire  _GEN_31; // @[IcmpNode.scala 247:26]
  wire  _GEN_32; // @[IcmpNode.scala 247:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UCMP FU ( // @[IcmpNode.scala 192:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[IcmpNode.scala 197:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[IcmpNode.scala 197:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[IcmpNode.scala 197:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[IcmpNode.scala 203:27]
  assign _GEN_12 = _T_117 ? 32'h8 : right_R_data; // @[IcmpNode.scala 203:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[IcmpNode.scala 203:27]
  assign _T_119 = left_R_taskID | right_R_taskID; // @[IcmpNode.scala 218:44]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[IcmpNode.scala 227:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[IcmpNode.scala 230:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[IcmpNode.scala 227:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[IcmpNode.scala 227:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[IcmpNode.scala 227:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[IcmpNode.scala 226:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[IcmpNode.scala 226:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[IcmpNode.scala 226:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[IcmpNode.scala 247:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[IcmpNode.scala 247:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[IcmpNode.scala 247:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[IcmpNode.scala 247:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[IcmpNode.scala 247:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_119 | enable_R_taskID; // @[IcmpNode.scala 217:20 IcmpNode.scala 218:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[IcmpNode.scala 217:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[IcmpNode.scala 196:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[IcmpNode.scala 202:20]
  assign FU_io_in1 = left_R_data; // @[IcmpNode.scala 193:13]
  assign FU_io_in2 = right_R_data; // @[IcmpNode.scala 194:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h8;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module CBranchNodeVariable(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [9:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output [9:0]  io_TrueOutput_0_bits_taskID,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [9:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [9:0] cmp_R_taskID; // @[BranchNode.scala 1295:22]
  reg [31:0] _RAND_0;
  reg  cmp_R_control; // @[BranchNode.scala 1295:22]
  reg [31:0] _RAND_1;
  reg  cmp_valid; // @[BranchNode.scala 1296:26]
  reg [31:0] _RAND_2;
  reg [9:0] enable_R_taskID; // @[BranchNode.scala 1299:25]
  reg [31:0] _RAND_3;
  reg  enable_R_control; // @[BranchNode.scala 1299:25]
  reg [31:0] _RAND_4;
  reg  enable_valid_R; // @[BranchNode.scala 1300:31]
  reg [31:0] _RAND_5;
  reg [9:0] output_true_R_taskID; // @[BranchNode.scala 1306:30]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1306:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1307:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1308:46]
  reg [31:0] _RAND_9;
  reg [9:0] output_false_R_taskID; // @[BranchNode.scala 1310:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1310:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1311:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1312:48]
  reg [31:0] _RAND_13;
  wire [9:0] task_id; // @[BranchNode.scala 1314:33]
  wire  _T_127; // @[Decoupled.scala 37:37]
  wire  _T_129; // @[BranchNode.scala 1320:44]
  wire  _GEN_1; // @[BranchNode.scala 1319:23]
  wire [9:0] _GEN_2; // @[BranchNode.scala 1319:23]
  wire  _GEN_3; // @[BranchNode.scala 1319:23]
  wire  _T_132; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_4; // @[BranchNode.scala 1345:24]
  wire  _GEN_5; // @[BranchNode.scala 1345:24]
  wire  _GEN_6; // @[BranchNode.scala 1345:24]
  wire  predicate; // @[BranchNode.scala 1351:36]
  wire  true_output; // @[BranchNode.scala 1352:31]
  wire  _T_134; // @[BranchNode.scala 1353:35]
  wire  false_output; // @[BranchNode.scala 1353:32]
  wire  _T_136; // @[Decoupled.scala 37:37]
  wire  _GEN_7; // @[BranchNode.scala 1366:33]
  wire  _GEN_8; // @[BranchNode.scala 1366:33]
  wire  _T_139; // @[Decoupled.scala 37:37]
  wire  _GEN_9; // @[BranchNode.scala 1384:34]
  wire  _GEN_10; // @[BranchNode.scala 1384:34]
  reg  state; // @[BranchNode.scala 1396:22]
  reg [31:0] _RAND_14;
  wire  _T_143; // @[Conditional.scala 37:30]
  wire  _T_144; // @[BranchNode.scala 1402:27]
  wire  _GEN_11; // @[BranchNode.scala 1402:65]
  wire  _GEN_12; // @[BranchNode.scala 1402:65]
  wire  _GEN_13; // @[BranchNode.scala 1402:65]
  wire  _T_151; // @[BranchNode.scala 1436:27]
  wire [9:0] _GEN_14; // @[BranchNode.scala 1436:47]
  wire  _GEN_15; // @[BranchNode.scala 1436:47]
  wire  _GEN_16; // @[BranchNode.scala 1436:47]
  wire  _GEN_17; // @[BranchNode.scala 1436:47]
  wire [9:0] _GEN_18; // @[BranchNode.scala 1436:47]
  wire  _GEN_19; // @[BranchNode.scala 1436:47]
  wire  _GEN_20; // @[BranchNode.scala 1436:47]
  wire [9:0] _GEN_21; // @[BranchNode.scala 1436:47]
  wire  _GEN_22; // @[BranchNode.scala 1436:47]
  wire  _GEN_23; // @[BranchNode.scala 1436:47]
  wire  _GEN_24; // @[BranchNode.scala 1436:47]
  wire  _GEN_26; // @[BranchNode.scala 1436:47]
  wire  _GEN_27; // @[BranchNode.scala 1436:47]
  wire  _GEN_28; // @[BranchNode.scala 1436:47]
  wire [9:0] _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_32; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_47; // @[Conditional.scala 40:58]
  wire  _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_49; // @[Conditional.scala 40:58]
  wire  _GEN_50; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire [9:0] _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  wire  _GEN_56; // @[Conditional.scala 40:58]
  wire  _GEN_58; // @[Conditional.scala 40:58]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1314:33]
  assign _T_127 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 37:37]
  assign _T_129 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1320:44]
  assign _GEN_1 = _T_127 ? _T_129 : cmp_R_control; // @[BranchNode.scala 1319:23]
  assign _GEN_2 = _T_127 ? io_CmpIO_bits_taskID : cmp_R_taskID; // @[BranchNode.scala 1319:23]
  assign _GEN_3 = _T_127 ? 1'h1 : cmp_valid; // @[BranchNode.scala 1319:23]
  assign _T_132 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_132 ? io_enable_bits_taskID : enable_R_taskID; // @[BranchNode.scala 1345:24]
  assign _GEN_5 = _T_132 ? io_enable_bits_control : enable_R_control; // @[BranchNode.scala 1345:24]
  assign _GEN_6 = _T_132 ? 1'h1 : enable_valid_R; // @[BranchNode.scala 1345:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1351:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1352:31]
  assign _T_134 = ~ cmp_R_control; // @[BranchNode.scala 1353:35]
  assign false_output = predicate & _T_134; // @[BranchNode.scala 1353:32]
  assign _T_136 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_136 ? 1'h1 : fire_true_R_0; // @[BranchNode.scala 1366:33]
  assign _GEN_8 = _T_136 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1366:33]
  assign _T_139 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_139 ? 1'h1 : fire_false_R_0; // @[BranchNode.scala 1384:34]
  assign _GEN_10 = _T_139 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1384:34]
  assign _T_143 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_144 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1402:27]
  assign _GEN_11 = _T_144 ? 1'h1 : _GEN_8; // @[BranchNode.scala 1402:65]
  assign _GEN_12 = _T_144 ? 1'h1 : _GEN_10; // @[BranchNode.scala 1402:65]
  assign _GEN_13 = _T_144 ? 1'h1 : state; // @[BranchNode.scala 1402:65]
  assign _T_151 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1436:27]
  assign _GEN_14 = _T_151 ? 10'h0 : _GEN_2; // @[BranchNode.scala 1436:47]
  assign _GEN_15 = _T_151 ? 1'h0 : _GEN_1; // @[BranchNode.scala 1436:47]
  assign _GEN_16 = _T_151 ? 1'h0 : _GEN_3; // @[BranchNode.scala 1436:47]
  assign _GEN_17 = _T_151 ? 1'h0 : _GEN_5; // @[BranchNode.scala 1436:47]
  assign _GEN_18 = _T_151 ? 10'h0 : _GEN_4; // @[BranchNode.scala 1436:47]
  assign _GEN_19 = _T_151 ? 1'h0 : _GEN_6; // @[BranchNode.scala 1436:47]
  assign _GEN_20 = _T_151 ? 1'h0 : true_output; // @[BranchNode.scala 1436:47]
  assign _GEN_21 = _T_151 ? 10'h0 : task_id; // @[BranchNode.scala 1436:47]
  assign _GEN_22 = _T_151 ? 1'h0 : _GEN_8; // @[BranchNode.scala 1436:47]
  assign _GEN_23 = _T_151 ? 1'h0 : _GEN_7; // @[BranchNode.scala 1436:47]
  assign _GEN_24 = _T_151 ? 1'h0 : false_output; // @[BranchNode.scala 1436:47]
  assign _GEN_26 = _T_151 ? 1'h0 : _GEN_10; // @[BranchNode.scala 1436:47]
  assign _GEN_27 = _T_151 ? 1'h0 : _GEN_9; // @[BranchNode.scala 1436:47]
  assign _GEN_28 = _T_151 ? 1'h0 : state; // @[BranchNode.scala 1436:47]
  assign _GEN_29 = state ? _GEN_14 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_30 = state ? _GEN_15 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_31 = state ? _GEN_16 : _GEN_3; // @[Conditional.scala 39:67]
  assign _GEN_32 = state ? _GEN_17 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_33 = state ? _GEN_18 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_19 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_20 : true_output; // @[Conditional.scala 39:67]
  assign _GEN_36 = state ? _GEN_21 : task_id; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_22 : _GEN_8; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_23 : _GEN_7; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_24 : false_output; // @[Conditional.scala 39:67]
  assign _GEN_41 = state ? _GEN_26 : _GEN_10; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_28 : state; // @[Conditional.scala 39:67]
  assign _GEN_44 = _T_143 ? _GEN_11 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_143 ? _GEN_12 : _GEN_41; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_143 ? _GEN_13 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_143 ? _GEN_2 : _GEN_29; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_143 ? _GEN_1 : _GEN_30; // @[Conditional.scala 40:58]
  assign _GEN_49 = _T_143 ? _GEN_3 : _GEN_31; // @[Conditional.scala 40:58]
  assign _GEN_50 = _T_143 ? _GEN_5 : _GEN_32; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_143 ? _GEN_4 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_143 ? _GEN_6 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_143 ? true_output : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_143 ? task_id : _GEN_36; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_143 ? _GEN_7 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_56 = _T_143 ? false_output : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_58 = _T_143 ? _GEN_9 : _GEN_42; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1344:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1318:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1362:28]
  assign io_TrueOutput_0_bits_taskID = output_true_R_taskID; // @[BranchNode.scala 1361:27]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1361:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1380:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1379:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1379:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_true_R_taskID = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cmp_R_taskID <= 10'h0;
    end else begin
      if (_T_143) begin
        if (_T_127) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            cmp_R_taskID <= 10'h0;
          end else begin
            if (_T_127) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_127) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_127) begin
          cmp_R_control <= _T_129;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_127) begin
              cmp_R_control <= _T_129;
            end
          end
        end else begin
          if (_T_127) begin
            cmp_R_control <= _T_129;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_127) begin
          cmp_valid <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            cmp_valid <= 1'h0;
          end else begin
            if (_T_127) begin
              cmp_valid <= 1'h1;
            end
          end
        end else begin
          if (_T_127) begin
            cmp_valid <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_143) begin
        if (_T_132) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            enable_R_taskID <= 10'h0;
          end else begin
            if (_T_132) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_132) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_132) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_132) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_132) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_132) begin
          enable_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_132) begin
              enable_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_132) begin
            enable_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_true_R_taskID <= 10'h0;
    end else begin
      if (_T_143) begin
        output_true_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_151) begin
            output_true_R_taskID <= 10'h0;
          end else begin
            output_true_R_taskID <= task_id;
          end
        end else begin
          output_true_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_143) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_151) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_144) begin
          output_true_valid_R_0 <= 1'h1;
        end else begin
          if (_T_136) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_136) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_136) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_136) begin
          fire_true_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            if (_T_136) begin
              fire_true_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_136) begin
            fire_true_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 10'h0;
    end else begin
      if (_T_143) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_151) begin
            output_false_R_taskID <= 10'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_143) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_151) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_144) begin
          output_false_valid_R_0 <= 1'h1;
        end else begin
          if (_T_139) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_139) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_139) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_139) begin
          fire_false_R_0 <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            if (_T_139) begin
              fire_false_R_0 <= 1'h1;
            end
          end
        end else begin
          if (_T_139) begin
            fire_false_R_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_143) begin
        if (_T_144) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_151) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_10(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_6;
  wire  _T_86; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 186:29]
  wire  _GEN_3; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_5; // @[HandShaking.scala 197:27]
  wire  _GEN_6; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_7;
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_9;
  reg [9:0] right_R_taskID; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_10;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_11;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_14;
  wire  _T_126; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_9; // @[ComputeNode.scala 77:26]
  wire [31:0] _GEN_10; // @[ComputeNode.scala 77:26]
  wire  _GEN_11; // @[ComputeNode.scala 77:26]
  wire  _T_129; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_13; // @[ComputeNode.scala 83:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 83:27]
  wire  _GEN_15; // @[ComputeNode.scala 83:27]
  wire [9:0] _T_131; // @[ComputeNode.scala 98:44]
  wire  _T_135; // @[Conditional.scala 37:30]
  wire  _T_136; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 110:34]
  wire  _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_20; // @[ComputeNode.scala 107:45]
  wire  _GEN_21; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_22; // @[ComputeNode.scala 107:45]
  wire  _GEN_25; // @[ComputeNode.scala 106:28]
  wire  _GEN_26; // @[ComputeNode.scala 106:28]
  wire  _GEN_27; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_28; // @[ComputeNode.scala 106:28]
  wire  _T_147; // @[HandShaking.scala 222:83]
  wire  _T_148; // @[HandShaking.scala 222:83]
  wire  _T_149; // @[HandShaking.scala 224:11]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[ComputeNode.scala 123:26]
  wire  _GEN_35; // @[ComputeNode.scala 123:26]
  wire  _GEN_36; // @[ComputeNode.scala 123:26]
  wire  _GEN_37; // @[ComputeNode.scala 123:26]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire  _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_86 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_86 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_86 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_88 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_88 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 186:29]
  assign _GEN_3 = _T_88 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_5 = _T_91 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_6 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_126 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_126 ? io_LeftIO_bits_taskID : left_R_taskID; // @[ComputeNode.scala 77:26]
  assign _GEN_10 = _T_126 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_11 = _T_126 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_129 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_13 = _T_129 ? io_RightIO_bits_taskID : right_R_taskID; // @[ComputeNode.scala 83:27]
  assign _GEN_14 = _T_129 ? 32'h1 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_15 = _T_129 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_131 = left_R_taskID | right_R_taskID; // @[ComputeNode.scala 98:44]
  assign _T_135 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_136 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_16 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_19 = _T_136 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_20 = _T_136 ? 1'h1 : _GEN_3; // @[ComputeNode.scala 107:45]
  assign _GEN_21 = _T_136 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = _T_136 ? _GEN_16 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_25 = enable_valid_R ? _GEN_19 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_26 = enable_valid_R ? _GEN_20 : _GEN_3; // @[ComputeNode.scala 106:28]
  assign _GEN_27 = enable_valid_R ? _GEN_21 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_28 = enable_valid_R ? _GEN_22 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_147 = out_ready_R_0 | _T_86; // @[HandShaking.scala 222:83]
  assign _T_148 = out_ready_R_1 | _T_88; // @[HandShaking.scala 222:83]
  assign _T_149 = _T_147 & _T_148; // @[HandShaking.scala 224:11]
  assign _GEN_31 = _T_149 ? 1'h0 : _GEN_11; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_149 ? 1'h0 : _GEN_15; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = _T_149 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_35 = _T_149 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_36 = _T_149 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_37 = _T_149 ? 1'h0 : _GEN_4; // @[ComputeNode.scala 123:26]
  assign _GEN_38 = state ? _GEN_31 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_32 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_33 : state; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_35 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_36 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_44 = state ? _GEN_37 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_45 = _T_135 ? _GEN_25 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_135 ? _GEN_26 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_135 ? _GEN_27 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_135 ? _GEN_28 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_135 ? _GEN_11 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_135 ? _GEN_15 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_135 ? _GEN_0 : _GEN_42; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_135 ? _GEN_2 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_135 ? _GEN_4 : _GEN_44; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 184:21]
  assign io_Out_1_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_1_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_R_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_valid_R = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_91) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_86) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_86) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_86) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_88) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_86) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_86) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_86) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_1 <= 1'h1;
          end else begin
            if (_T_88) begin
              out_valid_R_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_88) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_126) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_126) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_126) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_129) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_129) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_129) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_129) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_129) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module IcmpNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_in2; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_out; // @[IcmpNode.scala 192:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[IcmpNode.scala 170:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[IcmpNode.scala 174:30]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R_data; // @[IcmpNode.scala 179:27]
  reg [31:0] _RAND_11;
  reg  state; // @[IcmpNode.scala 182:22]
  reg [31:0] _RAND_12;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[IcmpNode.scala 197:26]
  wire [31:0] _GEN_8; // @[IcmpNode.scala 197:26]
  wire  _GEN_9; // @[IcmpNode.scala 197:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[IcmpNode.scala 203:27]
  wire [31:0] _GEN_12; // @[IcmpNode.scala 203:27]
  wire  _GEN_13; // @[IcmpNode.scala 203:27]
  wire [9:0] _T_119; // @[IcmpNode.scala 218:44]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[IcmpNode.scala 227:27]
  wire [31:0] _GEN_14; // @[IcmpNode.scala 230:34]
  wire  _GEN_17; // @[IcmpNode.scala 227:45]
  wire  _GEN_18; // @[IcmpNode.scala 227:45]
  wire [31:0] _GEN_19; // @[IcmpNode.scala 227:45]
  wire  _GEN_22; // @[IcmpNode.scala 226:28]
  wire  _GEN_23; // @[IcmpNode.scala 226:28]
  wire [31:0] _GEN_24; // @[IcmpNode.scala 226:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[IcmpNode.scala 247:26]
  wire  _GEN_28; // @[IcmpNode.scala 247:26]
  wire  _GEN_29; // @[IcmpNode.scala 247:26]
  wire  _GEN_31; // @[IcmpNode.scala 247:26]
  wire  _GEN_32; // @[IcmpNode.scala 247:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UCMP FU ( // @[IcmpNode.scala 192:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[IcmpNode.scala 197:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[IcmpNode.scala 197:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[IcmpNode.scala 197:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[IcmpNode.scala 203:27]
  assign _GEN_12 = _T_117 ? 32'h8 : right_R_data; // @[IcmpNode.scala 203:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[IcmpNode.scala 203:27]
  assign _T_119 = left_R_taskID | right_R_taskID; // @[IcmpNode.scala 218:44]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[IcmpNode.scala 227:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[IcmpNode.scala 230:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[IcmpNode.scala 227:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[IcmpNode.scala 227:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[IcmpNode.scala 227:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[IcmpNode.scala 226:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[IcmpNode.scala 226:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[IcmpNode.scala 226:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[IcmpNode.scala 247:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[IcmpNode.scala 247:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[IcmpNode.scala 247:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[IcmpNode.scala 247:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[IcmpNode.scala 247:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_119 | enable_R_taskID; // @[IcmpNode.scala 217:20 IcmpNode.scala 218:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[IcmpNode.scala 217:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[IcmpNode.scala 196:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[IcmpNode.scala 202:20]
  assign FU_io_in1 = left_R_data; // @[IcmpNode.scala 193:13]
  assign FU_io_in2 = right_R_data; // @[IcmpNode.scala 194:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h8;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_11(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_6;
  wire  _T_86; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 186:29]
  wire  _GEN_3; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_5; // @[HandShaking.scala 197:27]
  wire  _GEN_6; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_7;
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_9;
  reg [9:0] right_R_taskID; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_10;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_11;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_14;
  wire  _T_126; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_9; // @[ComputeNode.scala 77:26]
  wire [31:0] _GEN_10; // @[ComputeNode.scala 77:26]
  wire  _GEN_11; // @[ComputeNode.scala 77:26]
  wire  _T_129; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_13; // @[ComputeNode.scala 83:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 83:27]
  wire  _GEN_15; // @[ComputeNode.scala 83:27]
  wire [9:0] _T_131; // @[ComputeNode.scala 98:44]
  wire  _T_135; // @[Conditional.scala 37:30]
  wire  _T_136; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 110:34]
  wire  _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_20; // @[ComputeNode.scala 107:45]
  wire  _GEN_21; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_22; // @[ComputeNode.scala 107:45]
  wire  _GEN_25; // @[ComputeNode.scala 106:28]
  wire  _GEN_26; // @[ComputeNode.scala 106:28]
  wire  _GEN_27; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_28; // @[ComputeNode.scala 106:28]
  wire  _T_147; // @[HandShaking.scala 222:83]
  wire  _T_148; // @[HandShaking.scala 222:83]
  wire  _T_149; // @[HandShaking.scala 224:11]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[ComputeNode.scala 123:26]
  wire  _GEN_35; // @[ComputeNode.scala 123:26]
  wire  _GEN_36; // @[ComputeNode.scala 123:26]
  wire  _GEN_37; // @[ComputeNode.scala 123:26]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire  _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_86 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_86 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_86 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_88 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_88 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 186:29]
  assign _GEN_3 = _T_88 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_5 = _T_91 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_6 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_126 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_126 ? io_LeftIO_bits_taskID : left_R_taskID; // @[ComputeNode.scala 77:26]
  assign _GEN_10 = _T_126 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_11 = _T_126 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_129 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_13 = _T_129 ? io_RightIO_bits_taskID : right_R_taskID; // @[ComputeNode.scala 83:27]
  assign _GEN_14 = _T_129 ? 32'h1 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_15 = _T_129 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_131 = left_R_taskID | right_R_taskID; // @[ComputeNode.scala 98:44]
  assign _T_135 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_136 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_16 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_19 = _T_136 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_20 = _T_136 ? 1'h1 : _GEN_3; // @[ComputeNode.scala 107:45]
  assign _GEN_21 = _T_136 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = _T_136 ? _GEN_16 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_25 = enable_valid_R ? _GEN_19 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_26 = enable_valid_R ? _GEN_20 : _GEN_3; // @[ComputeNode.scala 106:28]
  assign _GEN_27 = enable_valid_R ? _GEN_21 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_28 = enable_valid_R ? _GEN_22 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_147 = out_ready_R_0 | _T_86; // @[HandShaking.scala 222:83]
  assign _T_148 = out_ready_R_1 | _T_88; // @[HandShaking.scala 222:83]
  assign _T_149 = _T_147 & _T_148; // @[HandShaking.scala 224:11]
  assign _GEN_31 = _T_149 ? 1'h0 : _GEN_11; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_149 ? 1'h0 : _GEN_15; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = _T_149 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_35 = _T_149 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_36 = _T_149 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_37 = _T_149 ? 1'h0 : _GEN_4; // @[ComputeNode.scala 123:26]
  assign _GEN_38 = state ? _GEN_31 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_32 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_33 : state; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_35 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_36 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_44 = state ? _GEN_37 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_45 = _T_135 ? _GEN_25 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_135 ? _GEN_26 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_135 ? _GEN_27 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_135 ? _GEN_28 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_135 ? _GEN_11 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_135 ? _GEN_15 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_135 ? _GEN_0 : _GEN_42; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_135 ? _GEN_2 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_135 ? _GEN_4 : _GEN_44; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 184:21]
  assign io_Out_1_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_1_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_R_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_valid_R = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_91) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_86) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_86) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_86) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_88) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_86) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_86) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_86) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_1 <= 1'h1;
          end else begin
            if (_T_88) begin
              out_valid_R_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_88) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_126) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_126) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_126) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_129) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_129) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_129) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_129) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_129) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module IcmpNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_in2; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_out; // @[IcmpNode.scala 192:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[IcmpNode.scala 170:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[IcmpNode.scala 174:30]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R_data; // @[IcmpNode.scala 179:27]
  reg [31:0] _RAND_11;
  reg  state; // @[IcmpNode.scala 182:22]
  reg [31:0] _RAND_12;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[IcmpNode.scala 197:26]
  wire [31:0] _GEN_8; // @[IcmpNode.scala 197:26]
  wire  _GEN_9; // @[IcmpNode.scala 197:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[IcmpNode.scala 203:27]
  wire [31:0] _GEN_12; // @[IcmpNode.scala 203:27]
  wire  _GEN_13; // @[IcmpNode.scala 203:27]
  wire [9:0] _T_119; // @[IcmpNode.scala 218:44]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[IcmpNode.scala 227:27]
  wire [31:0] _GEN_14; // @[IcmpNode.scala 230:34]
  wire  _GEN_17; // @[IcmpNode.scala 227:45]
  wire  _GEN_18; // @[IcmpNode.scala 227:45]
  wire [31:0] _GEN_19; // @[IcmpNode.scala 227:45]
  wire  _GEN_22; // @[IcmpNode.scala 226:28]
  wire  _GEN_23; // @[IcmpNode.scala 226:28]
  wire [31:0] _GEN_24; // @[IcmpNode.scala 226:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[IcmpNode.scala 247:26]
  wire  _GEN_28; // @[IcmpNode.scala 247:26]
  wire  _GEN_29; // @[IcmpNode.scala 247:26]
  wire  _GEN_31; // @[IcmpNode.scala 247:26]
  wire  _GEN_32; // @[IcmpNode.scala 247:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UCMP FU ( // @[IcmpNode.scala 192:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[IcmpNode.scala 197:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[IcmpNode.scala 197:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[IcmpNode.scala 197:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[IcmpNode.scala 203:27]
  assign _GEN_12 = _T_117 ? 32'h40 : right_R_data; // @[IcmpNode.scala 203:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[IcmpNode.scala 203:27]
  assign _T_119 = left_R_taskID | right_R_taskID; // @[IcmpNode.scala 218:44]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[IcmpNode.scala 227:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[IcmpNode.scala 230:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[IcmpNode.scala 227:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[IcmpNode.scala 227:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[IcmpNode.scala 227:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[IcmpNode.scala 226:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[IcmpNode.scala 226:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[IcmpNode.scala 226:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[IcmpNode.scala 247:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[IcmpNode.scala 247:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[IcmpNode.scala 247:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[IcmpNode.scala 247:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[IcmpNode.scala 247:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_119 | enable_R_taskID; // @[IcmpNode.scala 217:20 IcmpNode.scala 218:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[IcmpNode.scala 217:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[IcmpNode.scala 196:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[IcmpNode.scala 202:20]
  assign FU_io_in1 = left_R_data; // @[IcmpNode.scala 193:13]
  assign FU_io_in2 = right_R_data; // @[IcmpNode.scala 194:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h40;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_12(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_6;
  wire  _T_86; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 186:29]
  wire  _GEN_3; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_5; // @[HandShaking.scala 197:27]
  wire  _GEN_6; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_7;
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_9;
  reg [9:0] right_R_taskID; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_10;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_11;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_14;
  wire  _T_126; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_9; // @[ComputeNode.scala 77:26]
  wire [31:0] _GEN_10; // @[ComputeNode.scala 77:26]
  wire  _GEN_11; // @[ComputeNode.scala 77:26]
  wire  _T_129; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_13; // @[ComputeNode.scala 83:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 83:27]
  wire  _GEN_15; // @[ComputeNode.scala 83:27]
  wire [9:0] _T_131; // @[ComputeNode.scala 98:44]
  wire  _T_135; // @[Conditional.scala 37:30]
  wire  _T_136; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 110:34]
  wire  _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_20; // @[ComputeNode.scala 107:45]
  wire  _GEN_21; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_22; // @[ComputeNode.scala 107:45]
  wire  _GEN_25; // @[ComputeNode.scala 106:28]
  wire  _GEN_26; // @[ComputeNode.scala 106:28]
  wire  _GEN_27; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_28; // @[ComputeNode.scala 106:28]
  wire  _T_147; // @[HandShaking.scala 222:83]
  wire  _T_148; // @[HandShaking.scala 222:83]
  wire  _T_149; // @[HandShaking.scala 224:11]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[ComputeNode.scala 123:26]
  wire  _GEN_35; // @[ComputeNode.scala 123:26]
  wire  _GEN_36; // @[ComputeNode.scala 123:26]
  wire  _GEN_37; // @[ComputeNode.scala 123:26]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire  _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_86 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_86 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_86 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_88 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_88 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 186:29]
  assign _GEN_3 = _T_88 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_5 = _T_91 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_6 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_126 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_126 ? io_LeftIO_bits_taskID : left_R_taskID; // @[ComputeNode.scala 77:26]
  assign _GEN_10 = _T_126 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_11 = _T_126 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_129 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_13 = _T_129 ? io_RightIO_bits_taskID : right_R_taskID; // @[ComputeNode.scala 83:27]
  assign _GEN_14 = _T_129 ? 32'h8 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_15 = _T_129 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_131 = left_R_taskID | right_R_taskID; // @[ComputeNode.scala 98:44]
  assign _T_135 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_136 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_16 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_19 = _T_136 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_20 = _T_136 ? 1'h1 : _GEN_3; // @[ComputeNode.scala 107:45]
  assign _GEN_21 = _T_136 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = _T_136 ? _GEN_16 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_25 = enable_valid_R ? _GEN_19 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_26 = enable_valid_R ? _GEN_20 : _GEN_3; // @[ComputeNode.scala 106:28]
  assign _GEN_27 = enable_valid_R ? _GEN_21 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_28 = enable_valid_R ? _GEN_22 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_147 = out_ready_R_0 | _T_86; // @[HandShaking.scala 222:83]
  assign _T_148 = out_ready_R_1 | _T_88; // @[HandShaking.scala 222:83]
  assign _T_149 = _T_147 & _T_148; // @[HandShaking.scala 224:11]
  assign _GEN_31 = _T_149 ? 1'h0 : _GEN_11; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_149 ? 1'h0 : _GEN_15; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = _T_149 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_35 = _T_149 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_36 = _T_149 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_37 = _T_149 ? 1'h0 : _GEN_4; // @[ComputeNode.scala 123:26]
  assign _GEN_38 = state ? _GEN_31 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_32 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_33 : state; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_35 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_36 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_44 = state ? _GEN_37 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_45 = _T_135 ? _GEN_25 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_135 ? _GEN_26 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_135 ? _GEN_27 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_135 ? _GEN_28 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_135 ? _GEN_11 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_135 ? _GEN_15 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_135 ? _GEN_0 : _GEN_42; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_135 ? _GEN_2 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_135 ? _GEN_4 : _GEN_44; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 184:21]
  assign io_Out_1_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_1_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_R_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_valid_R = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_91) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_86) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_86) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_86) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_88) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_86) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_86) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_86) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_1 <= 1'h1;
          end else begin
            if (_T_88) begin
              out_valid_R_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_88) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_126) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_126) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_126) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_129) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_129) begin
        right_R_data <= 32'h8;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_129) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_129) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_129) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module UCMP_3(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire  _T_15; // @[Comparision.scala 85:33]
  assign _T_15 = io_in1 < io_in2; // @[Comparision.scala 85:33]
  assign io_out = {{31'd0}, _T_15}; // @[Comparision.scala 90:10]
endmodule
module IcmpNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_in2; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_out; // @[IcmpNode.scala 192:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[IcmpNode.scala 170:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[IcmpNode.scala 174:30]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R_data; // @[IcmpNode.scala 179:27]
  reg [31:0] _RAND_11;
  reg  state; // @[IcmpNode.scala 182:22]
  reg [31:0] _RAND_12;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[IcmpNode.scala 197:26]
  wire [31:0] _GEN_8; // @[IcmpNode.scala 197:26]
  wire  _GEN_9; // @[IcmpNode.scala 197:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[IcmpNode.scala 203:27]
  wire [31:0] _GEN_12; // @[IcmpNode.scala 203:27]
  wire  _GEN_13; // @[IcmpNode.scala 203:27]
  wire [9:0] _T_119; // @[IcmpNode.scala 218:44]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[IcmpNode.scala 227:27]
  wire [31:0] _GEN_14; // @[IcmpNode.scala 230:34]
  wire  _GEN_17; // @[IcmpNode.scala 227:45]
  wire  _GEN_18; // @[IcmpNode.scala 227:45]
  wire [31:0] _GEN_19; // @[IcmpNode.scala 227:45]
  wire  _GEN_22; // @[IcmpNode.scala 226:28]
  wire  _GEN_23; // @[IcmpNode.scala 226:28]
  wire [31:0] _GEN_24; // @[IcmpNode.scala 226:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[IcmpNode.scala 247:26]
  wire  _GEN_28; // @[IcmpNode.scala 247:26]
  wire  _GEN_29; // @[IcmpNode.scala 247:26]
  wire  _GEN_31; // @[IcmpNode.scala 247:26]
  wire  _GEN_32; // @[IcmpNode.scala 247:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UCMP_3 FU ( // @[IcmpNode.scala 192:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[IcmpNode.scala 197:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[IcmpNode.scala 197:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[IcmpNode.scala 197:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[IcmpNode.scala 203:27]
  assign _GEN_12 = _T_117 ? 32'h40 : right_R_data; // @[IcmpNode.scala 203:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[IcmpNode.scala 203:27]
  assign _T_119 = left_R_taskID | right_R_taskID; // @[IcmpNode.scala 218:44]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[IcmpNode.scala 227:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[IcmpNode.scala 230:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[IcmpNode.scala 227:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[IcmpNode.scala 227:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[IcmpNode.scala 227:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[IcmpNode.scala 226:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[IcmpNode.scala 226:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[IcmpNode.scala 226:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[IcmpNode.scala 247:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[IcmpNode.scala 247:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[IcmpNode.scala 247:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[IcmpNode.scala 247:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[IcmpNode.scala 247:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_119 | enable_R_taskID; // @[IcmpNode.scala 217:20 IcmpNode.scala 218:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[IcmpNode.scala 217:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[IcmpNode.scala 196:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[IcmpNode.scala 202:20]
  assign FU_io_in1 = left_R_data; // @[IcmpNode.scala 193:13]
  assign FU_io_in2 = right_R_data; // @[IcmpNode.scala 194:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h40;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ComputeNode_13(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [9:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 72:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 72:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_6;
  wire  _T_86; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_88; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 186:29]
  wire  _GEN_3; // @[HandShaking.scala 186:29]
  wire  _T_91; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_5; // @[HandShaking.scala 197:27]
  wire  _GEN_6; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_7;
  reg [31:0] left_R_data; // @[ComputeNode.scala 49:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 50:29]
  reg [31:0] _RAND_9;
  reg [9:0] right_R_taskID; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_10;
  reg [31:0] right_R_data; // @[ComputeNode.scala 53:24]
  reg [31:0] _RAND_11;
  reg  right_valid_R; // @[ComputeNode.scala 54:30]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R_data; // @[ComputeNode.scala 59:27]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 62:22]
  reg [31:0] _RAND_14;
  wire  _T_126; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_9; // @[ComputeNode.scala 77:26]
  wire [31:0] _GEN_10; // @[ComputeNode.scala 77:26]
  wire  _GEN_11; // @[ComputeNode.scala 77:26]
  wire  _T_129; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_13; // @[ComputeNode.scala 83:27]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 83:27]
  wire  _GEN_15; // @[ComputeNode.scala 83:27]
  wire [9:0] _T_131; // @[ComputeNode.scala 98:44]
  wire  _T_135; // @[Conditional.scala 37:30]
  wire  _T_136; // @[ComputeNode.scala 107:27]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 110:34]
  wire  _GEN_19; // @[ComputeNode.scala 107:45]
  wire  _GEN_20; // @[ComputeNode.scala 107:45]
  wire  _GEN_21; // @[ComputeNode.scala 107:45]
  wire [31:0] _GEN_22; // @[ComputeNode.scala 107:45]
  wire  _GEN_25; // @[ComputeNode.scala 106:28]
  wire  _GEN_26; // @[ComputeNode.scala 106:28]
  wire  _GEN_27; // @[ComputeNode.scala 106:28]
  wire [31:0] _GEN_28; // @[ComputeNode.scala 106:28]
  wire  _T_147; // @[HandShaking.scala 222:83]
  wire  _T_148; // @[HandShaking.scala 222:83]
  wire  _T_149; // @[HandShaking.scala 224:11]
  wire  _GEN_31; // @[ComputeNode.scala 123:26]
  wire  _GEN_32; // @[ComputeNode.scala 123:26]
  wire  _GEN_33; // @[ComputeNode.scala 123:26]
  wire  _GEN_35; // @[ComputeNode.scala 123:26]
  wire  _GEN_36; // @[ComputeNode.scala 123:26]
  wire  _GEN_37; // @[ComputeNode.scala 123:26]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_40; // @[Conditional.scala 39:67]
  wire  _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_43; // @[Conditional.scala 39:67]
  wire  _GEN_44; // @[Conditional.scala 39:67]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58]
  wire  _GEN_51; // @[Conditional.scala 40:58]
  wire  _GEN_52; // @[Conditional.scala 40:58]
  wire  _GEN_53; // @[Conditional.scala 40:58]
  wire  _GEN_54; // @[Conditional.scala 40:58]
  wire  _GEN_55; // @[Conditional.scala 40:58]
  UALU_1 FU ( // @[ComputeNode.scala 72:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_86 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_86 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_86 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_88 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_88 ? io_Out_1_ready : out_ready_R_1; // @[HandShaking.scala 186:29]
  assign _GEN_3 = _T_88 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 186:29]
  assign _T_91 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_91 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_5 = _T_91 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_6 = _T_91 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_126 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_9 = _T_126 ? io_LeftIO_bits_taskID : left_R_taskID; // @[ComputeNode.scala 77:26]
  assign _GEN_10 = _T_126 ? io_LeftIO_bits_data : left_R_data; // @[ComputeNode.scala 77:26]
  assign _GEN_11 = _T_126 ? 1'h1 : left_valid_R; // @[ComputeNode.scala 77:26]
  assign _T_129 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_13 = _T_129 ? io_RightIO_bits_taskID : right_R_taskID; // @[ComputeNode.scala 83:27]
  assign _GEN_14 = _T_129 ? 32'h8 : right_R_data; // @[ComputeNode.scala 83:27]
  assign _GEN_15 = _T_129 ? 1'h1 : right_valid_R; // @[ComputeNode.scala 83:27]
  assign _T_131 = left_R_taskID | right_R_taskID; // @[ComputeNode.scala 98:44]
  assign _T_135 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_136 = left_valid_R & right_valid_R; // @[ComputeNode.scala 107:27]
  assign _GEN_16 = enable_R_control ? FU_io_out : 32'h0; // @[ComputeNode.scala 110:34]
  assign _GEN_19 = _T_136 ? 1'h1 : _GEN_1; // @[ComputeNode.scala 107:45]
  assign _GEN_20 = _T_136 ? 1'h1 : _GEN_3; // @[ComputeNode.scala 107:45]
  assign _GEN_21 = _T_136 ? 1'h1 : state; // @[ComputeNode.scala 107:45]
  assign _GEN_22 = _T_136 ? _GEN_16 : out_data_R_data; // @[ComputeNode.scala 107:45]
  assign _GEN_25 = enable_valid_R ? _GEN_19 : _GEN_1; // @[ComputeNode.scala 106:28]
  assign _GEN_26 = enable_valid_R ? _GEN_20 : _GEN_3; // @[ComputeNode.scala 106:28]
  assign _GEN_27 = enable_valid_R ? _GEN_21 : state; // @[ComputeNode.scala 106:28]
  assign _GEN_28 = enable_valid_R ? _GEN_22 : out_data_R_data; // @[ComputeNode.scala 106:28]
  assign _T_147 = out_ready_R_0 | _T_86; // @[HandShaking.scala 222:83]
  assign _T_148 = out_ready_R_1 | _T_88; // @[HandShaking.scala 222:83]
  assign _T_149 = _T_147 & _T_148; // @[HandShaking.scala 224:11]
  assign _GEN_31 = _T_149 ? 1'h0 : _GEN_11; // @[ComputeNode.scala 123:26]
  assign _GEN_32 = _T_149 ? 1'h0 : _GEN_15; // @[ComputeNode.scala 123:26]
  assign _GEN_33 = _T_149 ? 1'h0 : state; // @[ComputeNode.scala 123:26]
  assign _GEN_35 = _T_149 ? 1'h0 : _GEN_0; // @[ComputeNode.scala 123:26]
  assign _GEN_36 = _T_149 ? 1'h0 : _GEN_2; // @[ComputeNode.scala 123:26]
  assign _GEN_37 = _T_149 ? 1'h0 : _GEN_4; // @[ComputeNode.scala 123:26]
  assign _GEN_38 = state ? _GEN_31 : _GEN_11; // @[Conditional.scala 39:67]
  assign _GEN_39 = state ? _GEN_32 : _GEN_15; // @[Conditional.scala 39:67]
  assign _GEN_40 = state ? _GEN_33 : state; // @[Conditional.scala 39:67]
  assign _GEN_42 = state ? _GEN_35 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_43 = state ? _GEN_36 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_44 = state ? _GEN_37 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_45 = _T_135 ? _GEN_25 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_135 ? _GEN_26 : _GEN_3; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_135 ? _GEN_27 : _GEN_40; // @[Conditional.scala 40:58]
  assign _GEN_48 = _T_135 ? _GEN_28 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_51 = _T_135 ? _GEN_11 : _GEN_38; // @[Conditional.scala 40:58]
  assign _GEN_52 = _T_135 ? _GEN_15 : _GEN_39; // @[Conditional.scala 40:58]
  assign _GEN_53 = _T_135 ? _GEN_0 : _GEN_42; // @[Conditional.scala 40:58]
  assign _GEN_54 = _T_135 ? _GEN_2 : _GEN_43; // @[Conditional.scala 40:58]
  assign _GEN_55 = _T_135 ? _GEN_4 : _GEN_44; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 184:21]
  assign io_Out_1_bits_taskID = _T_131 | enable_R_taskID; // @[ComputeNode.scala 97:20 ComputeNode.scala 98:27]
  assign io_Out_1_bits_data = out_data_R_data; // @[ComputeNode.scala 97:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 76:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 82:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 73:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 74:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_R_taskID = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_taskID = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_valid_R = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_91) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_91) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_91) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_91) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_91) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_86) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_86) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_86) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_88) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_86) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_86) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_86) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            out_valid_R_1 <= 1'h1;
          end else begin
            if (_T_88) begin
              out_valid_R_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_88) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_126) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_126) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_126) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_126) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_126) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_129) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_129) begin
        right_R_data <= 32'h8;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_135) begin
        if (_T_129) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_129) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_129) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_135) begin
        if (enable_valid_R) begin
          if (_T_136) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_149) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module IcmpNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [9:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [9:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [9:0]  io_LeftIO_bits_taskID,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [9:0]  io_RightIO_bits_taskID
);
  wire [31:0] FU_io_in1; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_in2; // @[IcmpNode.scala 192:18]
  wire [31:0] FU_io_out; // @[IcmpNode.scala 192:18]
  reg [9:0] enable_R_taskID; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 169:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 173:46]
  reg [31:0] _RAND_4;
  wire  _T_76; // @[Decoupled.scala 37:37]
  wire  _GEN_0; // @[HandShaking.scala 186:29]
  wire  _GEN_1; // @[HandShaking.scala 186:29]
  wire  _T_79; // @[Decoupled.scala 37:37]
  wire  _GEN_2; // @[HandShaking.scala 197:27]
  wire [9:0] _GEN_3; // @[HandShaking.scala 197:27]
  wire  _GEN_4; // @[HandShaking.scala 197:27]
  reg [9:0] left_R_taskID; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_5;
  reg [31:0] left_R_data; // @[IcmpNode.scala 169:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[IcmpNode.scala 170:29]
  reg [31:0] _RAND_7;
  reg [9:0] right_R_taskID; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_8;
  reg [31:0] right_R_data; // @[IcmpNode.scala 173:24]
  reg [31:0] _RAND_9;
  reg  right_valid_R; // @[IcmpNode.scala 174:30]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R_data; // @[IcmpNode.scala 179:27]
  reg [31:0] _RAND_11;
  reg  state; // @[IcmpNode.scala 182:22]
  reg [31:0] _RAND_12;
  wire  _T_114; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_7; // @[IcmpNode.scala 197:26]
  wire [31:0] _GEN_8; // @[IcmpNode.scala 197:26]
  wire  _GEN_9; // @[IcmpNode.scala 197:26]
  wire  _T_117; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_11; // @[IcmpNode.scala 203:27]
  wire [31:0] _GEN_12; // @[IcmpNode.scala 203:27]
  wire  _GEN_13; // @[IcmpNode.scala 203:27]
  wire [9:0] _T_119; // @[IcmpNode.scala 218:44]
  wire  _T_121; // @[Conditional.scala 37:30]
  wire  _T_122; // @[IcmpNode.scala 227:27]
  wire [31:0] _GEN_14; // @[IcmpNode.scala 230:34]
  wire  _GEN_17; // @[IcmpNode.scala 227:45]
  wire  _GEN_18; // @[IcmpNode.scala 227:45]
  wire [31:0] _GEN_19; // @[IcmpNode.scala 227:45]
  wire  _GEN_22; // @[IcmpNode.scala 226:28]
  wire  _GEN_23; // @[IcmpNode.scala 226:28]
  wire [31:0] _GEN_24; // @[IcmpNode.scala 226:28]
  wire  _T_131; // @[HandShaking.scala 222:83]
  wire  _GEN_27; // @[IcmpNode.scala 247:26]
  wire  _GEN_28; // @[IcmpNode.scala 247:26]
  wire  _GEN_29; // @[IcmpNode.scala 247:26]
  wire  _GEN_31; // @[IcmpNode.scala 247:26]
  wire  _GEN_32; // @[IcmpNode.scala 247:26]
  wire  _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_39; // @[Conditional.scala 40:58]
  wire  _GEN_40; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58]
  wire  _GEN_44; // @[Conditional.scala 40:58]
  wire  _GEN_45; // @[Conditional.scala 40:58]
  wire  _GEN_46; // @[Conditional.scala 40:58]
  wire  _GEN_47; // @[Conditional.scala 40:58]
  UCMP_3 FU ( // @[IcmpNode.scala 192:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_76 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 37:37]
  assign _GEN_0 = _T_76 ? io_Out_0_ready : out_ready_R_0; // @[HandShaking.scala 186:29]
  assign _GEN_1 = _T_76 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 186:29]
  assign _T_79 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_2 = _T_79 ? io_enable_valid : enable_valid_R; // @[HandShaking.scala 197:27]
  assign _GEN_3 = _T_79 ? io_enable_bits_taskID : enable_R_taskID; // @[HandShaking.scala 197:27]
  assign _GEN_4 = _T_79 ? io_enable_bits_control : enable_R_control; // @[HandShaking.scala 197:27]
  assign _T_114 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_7 = _T_114 ? io_LeftIO_bits_taskID : left_R_taskID; // @[IcmpNode.scala 197:26]
  assign _GEN_8 = _T_114 ? io_LeftIO_bits_data : left_R_data; // @[IcmpNode.scala 197:26]
  assign _GEN_9 = _T_114 ? 1'h1 : left_valid_R; // @[IcmpNode.scala 197:26]
  assign _T_117 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 37:37]
  assign _GEN_11 = _T_117 ? io_RightIO_bits_taskID : right_R_taskID; // @[IcmpNode.scala 203:27]
  assign _GEN_12 = _T_117 ? 32'h40 : right_R_data; // @[IcmpNode.scala 203:27]
  assign _GEN_13 = _T_117 ? 1'h1 : right_valid_R; // @[IcmpNode.scala 203:27]
  assign _T_119 = left_R_taskID | right_R_taskID; // @[IcmpNode.scala 218:44]
  assign _T_121 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_122 = left_valid_R & right_valid_R; // @[IcmpNode.scala 227:27]
  assign _GEN_14 = enable_R_control ? FU_io_out : 32'h0; // @[IcmpNode.scala 230:34]
  assign _GEN_17 = _T_122 ? 1'h1 : _GEN_1; // @[IcmpNode.scala 227:45]
  assign _GEN_18 = _T_122 ? 1'h1 : state; // @[IcmpNode.scala 227:45]
  assign _GEN_19 = _T_122 ? _GEN_14 : out_data_R_data; // @[IcmpNode.scala 227:45]
  assign _GEN_22 = enable_valid_R ? _GEN_17 : _GEN_1; // @[IcmpNode.scala 226:28]
  assign _GEN_23 = enable_valid_R ? _GEN_18 : state; // @[IcmpNode.scala 226:28]
  assign _GEN_24 = enable_valid_R ? _GEN_19 : out_data_R_data; // @[IcmpNode.scala 226:28]
  assign _T_131 = out_ready_R_0 | _T_76; // @[HandShaking.scala 222:83]
  assign _GEN_27 = _T_131 ? 1'h0 : _GEN_9; // @[IcmpNode.scala 247:26]
  assign _GEN_28 = _T_131 ? 1'h0 : _GEN_13; // @[IcmpNode.scala 247:26]
  assign _GEN_29 = _T_131 ? 1'h0 : state; // @[IcmpNode.scala 247:26]
  assign _GEN_31 = _T_131 ? 1'h0 : _GEN_0; // @[IcmpNode.scala 247:26]
  assign _GEN_32 = _T_131 ? 1'h0 : _GEN_2; // @[IcmpNode.scala 247:26]
  assign _GEN_33 = state ? _GEN_27 : _GEN_9; // @[Conditional.scala 39:67]
  assign _GEN_34 = state ? _GEN_28 : _GEN_13; // @[Conditional.scala 39:67]
  assign _GEN_35 = state ? _GEN_29 : state; // @[Conditional.scala 39:67]
  assign _GEN_37 = state ? _GEN_31 : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_38 = state ? _GEN_32 : _GEN_2; // @[Conditional.scala 39:67]
  assign _GEN_39 = _T_121 ? _GEN_22 : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_40 = _T_121 ? _GEN_23 : _GEN_35; // @[Conditional.scala 40:58]
  assign _GEN_41 = _T_121 ? _GEN_24 : out_data_R_data; // @[Conditional.scala 40:58]
  assign _GEN_44 = _T_121 ? _GEN_9 : _GEN_33; // @[Conditional.scala 40:58]
  assign _GEN_45 = _T_121 ? _GEN_13 : _GEN_34; // @[Conditional.scala 40:58]
  assign _GEN_46 = _T_121 ? _GEN_0 : _GEN_37; // @[Conditional.scala 40:58]
  assign _GEN_47 = _T_121 ? _GEN_2 : _GEN_38; // @[Conditional.scala 40:58]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 196:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 184:21]
  assign io_Out_0_bits_taskID = _T_119 | enable_R_taskID; // @[IcmpNode.scala 217:20 IcmpNode.scala 218:27]
  assign io_Out_0_bits_data = out_data_R_data; // @[IcmpNode.scala 217:20]
  assign io_LeftIO_ready = ~ left_valid_R; // @[IcmpNode.scala 196:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[IcmpNode.scala 202:20]
  assign FU_io_in1 = left_R_data; // @[IcmpNode.scala 193:13]
  assign FU_io_in2 = right_R_data; // @[IcmpNode.scala 194:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  left_R_taskID = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_taskID = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_R_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_79) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_79) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_79) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_79) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_76) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            out_valid_R_0 <= 1'h1;
          end else begin
            if (_T_76) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_76) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      left_R_taskID <= 10'h0;
    end else begin
      if (_T_114) begin
        left_R_taskID <= io_LeftIO_bits_taskID;
      end
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_114) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_114) begin
          left_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            left_valid_R <= 1'h0;
          end else begin
            if (_T_114) begin
              left_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_114) begin
            left_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      right_R_taskID <= 10'h0;
    end else begin
      if (_T_117) begin
        right_R_taskID <= io_RightIO_bits_taskID;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_117) begin
        right_R_data <= 32'h40;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_121) begin
        if (_T_117) begin
          right_valid_R <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            right_valid_R <= 1'h0;
          end else begin
            if (_T_117) begin
              right_valid_R <= 1'h1;
            end
          end
        end else begin
          if (_T_117) begin
            right_valid_R <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      out_data_R_data <= 32'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            if (enable_R_control) begin
              out_data_R_data <= FU_io_out;
            end else begin
              out_data_R_data <= 32'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_121) begin
        if (enable_valid_R) begin
          if (_T_122) begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_131) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module RetNode2(
  input        clock,
  input        reset,
  output       io_In_enable_ready,
  input        io_In_enable_valid,
  input  [9:0] io_In_enable_bits_taskID,
  input        io_In_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid,
  output [9:0] io_Out_bits_enable_taskID,
  output       io_Out_bits_enable_control
);
  reg  state; // @[RetNode.scala 236:22]
  reg [31:0] _RAND_0;
  reg  enable_valid_R; // @[RetNode.scala 239:31]
  reg [31:0] _RAND_1;
  reg [9:0] output_R_enable_taskID; // @[RetNode.scala 245:25]
  reg [31:0] _RAND_2;
  reg  output_R_enable_control; // @[RetNode.scala 245:25]
  reg [31:0] _RAND_3;
  reg  out_ready_R; // @[RetNode.scala 246:28]
  reg [31:0] _RAND_4;
  reg  out_valid_R; // @[RetNode.scala 247:28]
  reg [31:0] _RAND_5;
  wire  _T_39; // @[Decoupled.scala 37:37]
  wire  _GEN_1; // @[RetNode.scala 259:29]
  wire  _GEN_2; // @[RetNode.scala 259:29]
  wire [9:0] _GEN_3; // @[RetNode.scala 259:29]
  wire  _T_40; // @[Decoupled.scala 37:37]
  wire  _GEN_4; // @[RetNode.scala 277:23]
  wire  _GEN_5; // @[RetNode.scala 277:23]
  wire  _T_42; // @[Conditional.scala 37:30]
  wire  _GEN_8; // @[RetNode.scala 284:28]
  wire  _GEN_9; // @[RetNode.scala 284:28]
  wire  _GEN_10; // @[RetNode.scala 292:25]
  wire  _GEN_11; // @[RetNode.scala 292:25]
  wire  _GEN_12; // @[RetNode.scala 292:25]
  wire  _GEN_13; // @[RetNode.scala 292:25]
  wire  _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_16; // @[Conditional.scala 39:67]
  wire  _GEN_17; // @[Conditional.scala 39:67]
  wire  _GEN_18; // @[Conditional.scala 40:58]
  wire  _GEN_19; // @[Conditional.scala 40:58]
  wire  _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_21; // @[Conditional.scala 40:58]
  assign _T_39 = io_In_enable_ready & io_In_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_1 = _T_39 ? io_In_enable_valid : enable_valid_R; // @[RetNode.scala 259:29]
  assign _GEN_2 = _T_39 ? io_In_enable_bits_control : output_R_enable_control; // @[RetNode.scala 259:29]
  assign _GEN_3 = _T_39 ? io_In_enable_bits_taskID : output_R_enable_taskID; // @[RetNode.scala 259:29]
  assign _T_40 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 37:37]
  assign _GEN_4 = _T_40 ? io_Out_ready : out_ready_R; // @[RetNode.scala 277:23]
  assign _GEN_5 = _T_40 ? 1'h0 : out_valid_R; // @[RetNode.scala 277:23]
  assign _T_42 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_8 = enable_valid_R ? 1'h1 : _GEN_5; // @[RetNode.scala 284:28]
  assign _GEN_9 = enable_valid_R ? 1'h1 : state; // @[RetNode.scala 284:28]
  assign _GEN_10 = out_ready_R ? 1'h0 : _GEN_5; // @[RetNode.scala 292:25]
  assign _GEN_11 = out_ready_R ? 1'h0 : _GEN_1; // @[RetNode.scala 292:25]
  assign _GEN_12 = out_ready_R ? 1'h0 : _GEN_4; // @[RetNode.scala 292:25]
  assign _GEN_13 = out_ready_R ? 1'h0 : state; // @[RetNode.scala 292:25]
  assign _GEN_14 = state ? _GEN_10 : _GEN_5; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_11 : _GEN_1; // @[Conditional.scala 39:67]
  assign _GEN_16 = state ? _GEN_12 : _GEN_4; // @[Conditional.scala 39:67]
  assign _GEN_17 = state ? _GEN_13 : state; // @[Conditional.scala 39:67]
  assign _GEN_18 = _T_42 ? _GEN_8 : _GEN_14; // @[Conditional.scala 40:58]
  assign _GEN_19 = _T_42 ? _GEN_9 : _GEN_17; // @[Conditional.scala 40:58]
  assign _GEN_20 = _T_42 ? _GEN_1 : _GEN_15; // @[Conditional.scala 40:58]
  assign _GEN_21 = _T_42 ? _GEN_4 : _GEN_16; // @[Conditional.scala 40:58]
  assign io_In_enable_ready = ~ enable_valid_R; // @[RetNode.scala 258:22]
  assign io_Out_valid = out_valid_R; // @[RetNode.scala 275:16]
  assign io_Out_bits_enable_taskID = output_R_enable_taskID; // @[RetNode.scala 274:15]
  assign io_Out_bits_enable_control = output_R_enable_control; // @[RetNode.scala 274:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_valid_R = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  output_R_enable_taskID = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  output_R_enable_control = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_42) begin
        if (enable_valid_R) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_42) begin
        if (_T_39) begin
          enable_valid_R <= io_In_enable_valid;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_39) begin
              enable_valid_R <= io_In_enable_valid;
            end
          end
        end else begin
          if (_T_39) begin
            enable_valid_R <= io_In_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      output_R_enable_taskID <= 10'h0;
    end else begin
      if (_T_39) begin
        output_R_enable_taskID <= io_In_enable_bits_taskID;
      end
    end
    if (reset) begin
      output_R_enable_control <= 1'h0;
    end else begin
      if (_T_39) begin
        output_R_enable_control <= io_In_enable_bits_control;
      end
    end
    if (reset) begin
      out_ready_R <= 1'h0;
    end else begin
      if (_T_42) begin
        if (_T_40) begin
          out_ready_R <= io_Out_ready;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            out_ready_R <= 1'h0;
          end else begin
            if (_T_40) begin
              out_ready_R <= io_Out_ready;
            end
          end
        end else begin
          if (_T_40) begin
            out_ready_R <= io_Out_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R <= 1'h0;
    end else begin
      if (_T_42) begin
        if (enable_valid_R) begin
          out_valid_R <= 1'h1;
        end else begin
          if (_T_40) begin
            out_valid_R <= 1'h0;
          end
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            out_valid_R <= 1'h0;
          end else begin
            if (_T_40) begin
              out_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_40) begin
            out_valid_R <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ConstFastNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [9:0] io_Out_bits_taskID
);
  reg [9:0] enable_R_taskID; // @[ConstNode.scala 109:25]
  reg [31:0] _RAND_0;
  wire [9:0] task_input; // @[ConstNode.scala 112:43]
  reg  state; // @[ConstNode.scala 133:22]
  reg [31:0] _RAND_1;
  wire  _T_43; // @[Conditional.scala 37:30]
  wire  _T_46; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[ConstNode.scala 140:30]
  wire [9:0] _GEN_4; // @[ConstNode.scala 140:30]
  wire  _GEN_6; // @[ConstNode.scala 140:30]
  wire  _T_50; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_8; // @[ConstNode.scala 160:25]
  wire  _GEN_10; // @[ConstNode.scala 160:25]
  wire [9:0] _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ConstNode.scala 112:43]
  assign _T_43 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_46 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_46 ? io_enable_bits_taskID : task_input; // @[ConstNode.scala 140:30]
  assign _GEN_4 = _T_46 ? io_enable_bits_taskID : enable_R_taskID; // @[ConstNode.scala 140:30]
  assign _GEN_6 = _T_46 ? 1'h1 : state; // @[ConstNode.scala 140:30]
  assign _T_50 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_50 ? 10'h0 : enable_R_taskID; // @[ConstNode.scala 160:25]
  assign _GEN_10 = _T_50 ? 1'h0 : state; // @[ConstNode.scala 160:25]
  assign _GEN_13 = state ? _GEN_8 : enable_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : state; // @[Conditional.scala 39:67]
  assign _GEN_20 = _T_43 ? _GEN_4 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_43 ? _GEN_6 : _GEN_15; // @[Conditional.scala 40:58]
  assign io_enable_ready = 1'h0 == state; // @[ConstNode.scala 122:19 ConstNode.scala 137:23]
  assign io_Out_valid = _T_43 ? _T_46 : state; // @[ConstNode.scala 127:16 ConstNode.scala 138:20 ConstNode.scala 142:22 ConstNode.scala 158:20]
  assign io_Out_bits_taskID = _T_43 ? _GEN_3 : task_input; // @[ConstNode.scala 126:22 ConstNode.scala 144:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            enable_R_taskID <= 10'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ConstFastNode_3(
  input   clock,
  input   reset,
  output  io_enable_ready,
  input   io_enable_valid,
  input   io_Out_ready,
  output  io_Out_valid
);
  reg  state; // @[ConstNode.scala 133:22]
  reg [31:0] _RAND_0;
  wire  _T_43; // @[Conditional.scala 37:30]
  wire  _T_46; // @[Decoupled.scala 37:37]
  wire  _GEN_6; // @[ConstNode.scala 140:30]
  wire  _T_50; // @[Decoupled.scala 37:37]
  wire  _GEN_10; // @[ConstNode.scala 160:25]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  assign _T_43 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_46 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_6 = _T_46 ? 1'h1 : state; // @[ConstNode.scala 140:30]
  assign _T_50 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 37:37]
  assign _GEN_10 = _T_50 ? 1'h0 : state; // @[ConstNode.scala 160:25]
  assign _GEN_15 = state ? _GEN_10 : state; // @[Conditional.scala 39:67]
  assign _GEN_22 = _T_43 ? _GEN_6 : _GEN_15; // @[Conditional.scala 40:58]
  assign io_enable_ready = 1'h0 == state; // @[ConstNode.scala 122:19 ConstNode.scala 137:23]
  assign io_Out_valid = _T_43 ? _T_46 : state; // @[ConstNode.scala 127:16 ConstNode.scala 138:20 ConstNode.scala 142:22 ConstNode.scala 158:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ConstFastNode_7(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [9:0] io_Out_bits_taskID
);
  reg [9:0] enable_R_taskID; // @[ConstNode.scala 109:25]
  reg [31:0] _RAND_0;
  wire [9:0] task_input; // @[ConstNode.scala 112:43]
  reg  state; // @[ConstNode.scala 133:22]
  reg [31:0] _RAND_1;
  wire  _T_43; // @[Conditional.scala 37:30]
  wire  _T_46; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[ConstNode.scala 140:30]
  wire [9:0] _GEN_4; // @[ConstNode.scala 140:30]
  wire  _GEN_6; // @[ConstNode.scala 140:30]
  wire  _T_50; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_8; // @[ConstNode.scala 160:25]
  wire  _GEN_10; // @[ConstNode.scala 160:25]
  wire [9:0] _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ConstNode.scala 112:43]
  assign _T_43 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_46 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_46 ? io_enable_bits_taskID : task_input; // @[ConstNode.scala 140:30]
  assign _GEN_4 = _T_46 ? io_enable_bits_taskID : enable_R_taskID; // @[ConstNode.scala 140:30]
  assign _GEN_6 = _T_46 ? 1'h1 : state; // @[ConstNode.scala 140:30]
  assign _T_50 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_50 ? 10'h0 : enable_R_taskID; // @[ConstNode.scala 160:25]
  assign _GEN_10 = _T_50 ? 1'h0 : state; // @[ConstNode.scala 160:25]
  assign _GEN_13 = state ? _GEN_8 : enable_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : state; // @[Conditional.scala 39:67]
  assign _GEN_20 = _T_43 ? _GEN_4 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_43 ? _GEN_6 : _GEN_15; // @[Conditional.scala 40:58]
  assign io_enable_ready = 1'h0 == state; // @[ConstNode.scala 122:19 ConstNode.scala 137:23]
  assign io_Out_valid = _T_43 ? _T_46 : state; // @[ConstNode.scala 127:16 ConstNode.scala 138:20 ConstNode.scala 142:22 ConstNode.scala 158:20]
  assign io_Out_bits_taskID = _T_43 ? _GEN_3 : task_input; // @[ConstNode.scala 126:22 ConstNode.scala 144:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            enable_R_taskID <= 10'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ConstFastNode_8(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [9:0] io_Out_bits_taskID
);
  reg [9:0] enable_R_taskID; // @[ConstNode.scala 109:25]
  reg [31:0] _RAND_0;
  wire [9:0] task_input; // @[ConstNode.scala 112:43]
  reg  state; // @[ConstNode.scala 133:22]
  reg [31:0] _RAND_1;
  wire  _T_43; // @[Conditional.scala 37:30]
  wire  _T_46; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[ConstNode.scala 140:30]
  wire [9:0] _GEN_4; // @[ConstNode.scala 140:30]
  wire  _GEN_6; // @[ConstNode.scala 140:30]
  wire  _T_50; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_8; // @[ConstNode.scala 160:25]
  wire  _GEN_10; // @[ConstNode.scala 160:25]
  wire [9:0] _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ConstNode.scala 112:43]
  assign _T_43 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_46 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_46 ? io_enable_bits_taskID : task_input; // @[ConstNode.scala 140:30]
  assign _GEN_4 = _T_46 ? io_enable_bits_taskID : enable_R_taskID; // @[ConstNode.scala 140:30]
  assign _GEN_6 = _T_46 ? 1'h1 : state; // @[ConstNode.scala 140:30]
  assign _T_50 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_50 ? 10'h0 : enable_R_taskID; // @[ConstNode.scala 160:25]
  assign _GEN_10 = _T_50 ? 1'h0 : state; // @[ConstNode.scala 160:25]
  assign _GEN_13 = state ? _GEN_8 : enable_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : state; // @[Conditional.scala 39:67]
  assign _GEN_20 = _T_43 ? _GEN_4 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_43 ? _GEN_6 : _GEN_15; // @[Conditional.scala 40:58]
  assign io_enable_ready = 1'h0 == state; // @[ConstNode.scala 122:19 ConstNode.scala 137:23]
  assign io_Out_valid = _T_43 ? _T_46 : state; // @[ConstNode.scala 127:16 ConstNode.scala 138:20 ConstNode.scala 142:22 ConstNode.scala 158:20]
  assign io_Out_bits_taskID = _T_43 ? _GEN_3 : task_input; // @[ConstNode.scala 126:22 ConstNode.scala 144:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            enable_R_taskID <= 10'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module ConstFastNode_12(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [9:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [9:0] io_Out_bits_taskID
);
  reg [9:0] enable_R_taskID; // @[ConstNode.scala 109:25]
  reg [31:0] _RAND_0;
  wire [9:0] task_input; // @[ConstNode.scala 112:43]
  reg  state; // @[ConstNode.scala 133:22]
  reg [31:0] _RAND_1;
  wire  _T_43; // @[Conditional.scala 37:30]
  wire  _T_46; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_3; // @[ConstNode.scala 140:30]
  wire [9:0] _GEN_4; // @[ConstNode.scala 140:30]
  wire  _GEN_6; // @[ConstNode.scala 140:30]
  wire  _T_50; // @[Decoupled.scala 37:37]
  wire [9:0] _GEN_8; // @[ConstNode.scala 160:25]
  wire  _GEN_10; // @[ConstNode.scala 160:25]
  wire [9:0] _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_15; // @[Conditional.scala 39:67]
  wire [9:0] _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_22; // @[Conditional.scala 40:58]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ConstNode.scala 112:43]
  assign _T_43 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_46 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 37:37]
  assign _GEN_3 = _T_46 ? io_enable_bits_taskID : task_input; // @[ConstNode.scala 140:30]
  assign _GEN_4 = _T_46 ? io_enable_bits_taskID : enable_R_taskID; // @[ConstNode.scala 140:30]
  assign _GEN_6 = _T_46 ? 1'h1 : state; // @[ConstNode.scala 140:30]
  assign _T_50 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 37:37]
  assign _GEN_8 = _T_50 ? 10'h0 : enable_R_taskID; // @[ConstNode.scala 160:25]
  assign _GEN_10 = _T_50 ? 1'h0 : state; // @[ConstNode.scala 160:25]
  assign _GEN_13 = state ? _GEN_8 : enable_R_taskID; // @[Conditional.scala 39:67]
  assign _GEN_15 = state ? _GEN_10 : state; // @[Conditional.scala 39:67]
  assign _GEN_20 = _T_43 ? _GEN_4 : _GEN_13; // @[Conditional.scala 40:58]
  assign _GEN_22 = _T_43 ? _GEN_6 : _GEN_15; // @[Conditional.scala 40:58]
  assign io_enable_ready = 1'h0 == state; // @[ConstNode.scala 122:19 ConstNode.scala 137:23]
  assign io_Out_valid = _T_43 ? _T_46 : state; // @[ConstNode.scala 127:16 ConstNode.scala 138:20 ConstNode.scala 142:22 ConstNode.scala 158:20]
  assign io_Out_bits_taskID = _T_43 ? _GEN_3 : task_input; // @[ConstNode.scala 126:22 ConstNode.scala 144:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 10'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            enable_R_taskID <= 10'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          state <= 1'h1;
        end
      end else begin
        if (state) begin
          if (_T_50) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module bbgemmTop(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [9:0]  io_in_bits_enable_taskID,
  input         io_in_bits_enable_control,
  input         io_in_bits_data_field2_predicate,
  input  [9:0]  io_in_bits_data_field2_taskID,
  input  [31:0] io_in_bits_data_field2_data,
  input         io_in_bits_data_field1_predicate,
  input  [9:0]  io_in_bits_data_field1_taskID,
  input  [31:0] io_in_bits_data_field1_data,
  input         io_in_bits_data_field0_predicate,
  input  [9:0]  io_in_bits_data_field0_taskID,
  input  [31:0] io_in_bits_data_field0_data,
  input         io_MemResp_valid,
  input         io_MemResp_bits_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  input  [31:0] io_MemResp_bits_tile,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [9:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  output [31:0] io_MemReq_bits_tile,
  input         io_out_ready,
  output        io_out_valid,
  output [9:0]  io_out_bits_enable_taskID,
  output        io_out_bits_enable_control
);
  wire  MemCtrl_clock; // @[bbgemm.scala 45:23]
  wire  MemCtrl_reset; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_WriteIn_0_ready; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_WriteIn_0_valid; // @[bbgemm.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_0_bits_address; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_0_bits_data; // @[bbgemm.scala 45:23]
  wire [9:0] MemCtrl_io_WriteIn_0_bits_taskID; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_WriteOut_0_valid; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadIn_0_ready; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadIn_0_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_0_bits_address; // @[bbgemm.scala 45:23]
  wire [9:0] MemCtrl_io_ReadIn_0_bits_taskID; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadIn_1_ready; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadIn_1_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_1_bits_address; // @[bbgemm.scala 45:23]
  wire [9:0] MemCtrl_io_ReadIn_1_bits_taskID; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadIn_2_ready; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadIn_2_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_2_bits_address; // @[bbgemm.scala 45:23]
  wire [9:0] MemCtrl_io_ReadIn_2_bits_taskID; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadOut_0_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_0_data; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadOut_1_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_1_data; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_ReadOut_2_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_2_data; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_MemResp_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_MemResp_bits_data; // @[bbgemm.scala 45:23]
  wire [7:0] MemCtrl_io_MemResp_bits_tag; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_MemResp_bits_iswrite; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_MemReq_ready; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_MemReq_valid; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_MemReq_bits_addr; // @[bbgemm.scala 45:23]
  wire [31:0] MemCtrl_io_MemReq_bits_data; // @[bbgemm.scala 45:23]
  wire [3:0] MemCtrl_io_MemReq_bits_mask; // @[bbgemm.scala 45:23]
  wire [7:0] MemCtrl_io_MemReq_bits_tag; // @[bbgemm.scala 45:23]
  wire [9:0] MemCtrl_io_MemReq_bits_taskID; // @[bbgemm.scala 45:23]
  wire  MemCtrl_io_MemReq_bits_iswrite; // @[bbgemm.scala 45:23]
  wire  InputSplitter_clock; // @[bbgemm.scala 53:29]
  wire  InputSplitter_reset; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_In_ready; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_In_valid; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_In_bits_enable_taskID; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_In_bits_enable_control; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_In_bits_data_field2_taskID; // @[bbgemm.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field2_data; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_In_bits_data_field1_taskID; // @[bbgemm.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field1_data; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_In_bits_data_field0_taskID; // @[bbgemm.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field0_data; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_enable_ready; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_enable_valid; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_Out_enable_bits_taskID; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_enable_bits_control; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_data_field2_0_ready; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_data_field2_0_valid; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_Out_data_field2_0_bits_taskID; // @[bbgemm.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field2_0_bits_data; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_ready; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_valid; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_Out_data_field1_0_bits_taskID; // @[bbgemm.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_0_bits_data; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_data_field0_0_ready; // @[bbgemm.scala 53:29]
  wire  InputSplitter_io_Out_data_field0_0_valid; // @[bbgemm.scala 53:29]
  wire [9:0] InputSplitter_io_Out_data_field0_0_bits_taskID; // @[bbgemm.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field0_0_bits_data; // @[bbgemm.scala 53:29]
  wire  Loop_0_clock; // @[bbgemm.scala 62:22]
  wire  Loop_0_reset; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_enable_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_enable_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_enable_bits_taskID; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_enable_bits_control; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_0_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_1_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_1_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_InLiveIn_1_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_1_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_2_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_2_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_2_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_3_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_3_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_InLiveIn_3_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_3_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_4_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_4_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_InLiveIn_4_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_4_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_5_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_InLiveIn_5_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_5_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field5_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field5_1_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field5_1_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field5_1_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field4_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_OutLiveIn_field4_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_OutLiveIn_field3_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_activate_loop_start_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_activate_loop_start_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_activate_loop_start_bits_control; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_activate_loop_back_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_activate_loop_back_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_activate_loop_back_bits_control; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopBack_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopBack_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_loopBack_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopBack_0_bits_control; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopFinish_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopFinish_0_valid; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopFinish_0_bits_control; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopExit_0_ready; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopExit_0_valid; // @[bbgemm.scala 62:22]
  wire [9:0] Loop_0_io_loopExit_0_bits_taskID; // @[bbgemm.scala 62:22]
  wire  Loop_0_io_loopExit_0_bits_control; // @[bbgemm.scala 62:22]
  wire  Loop_1_clock; // @[bbgemm.scala 64:22]
  wire  Loop_1_reset; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_enable_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_enable_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_enable_bits_taskID; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_enable_bits_control; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_0_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_1_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_1_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_InLiveIn_1_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_1_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_2_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_2_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_InLiveIn_2_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_2_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_3_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_4_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_4_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_4_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_5_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_InLiveIn_5_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_InLiveIn_5_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_5_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field5_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_OutLiveIn_field5_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field4_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field4_1_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field4_1_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field4_1_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_1_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_1_valid; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field0_1_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_activate_loop_start_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_activate_loop_start_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_activate_loop_start_bits_control; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_activate_loop_back_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_activate_loop_back_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_activate_loop_back_bits_control; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopBack_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopBack_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_loopBack_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopBack_0_bits_control; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopFinish_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopFinish_0_valid; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopFinish_0_bits_control; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopExit_0_ready; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopExit_0_valid; // @[bbgemm.scala 64:22]
  wire [9:0] Loop_1_io_loopExit_0_bits_taskID; // @[bbgemm.scala 64:22]
  wire  Loop_1_io_loopExit_0_bits_control; // @[bbgemm.scala 64:22]
  wire  Loop_2_clock; // @[bbgemm.scala 66:22]
  wire  Loop_2_reset; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_enable_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_enable_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_enable_bits_taskID; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_enable_bits_control; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_0_valid; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_1_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_1_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_InLiveIn_1_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_1_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_2_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_2_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_InLiveIn_2_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_2_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_3_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_3_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_InLiveIn_3_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_3_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_4_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_InLiveIn_4_valid; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_4_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field4_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_OutLiveIn_field3_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_activate_loop_start_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_activate_loop_start_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_activate_loop_start_bits_control; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_activate_loop_back_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_activate_loop_back_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_activate_loop_back_bits_control; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopBack_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopBack_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_loopBack_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopBack_0_bits_control; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopFinish_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopFinish_0_valid; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopFinish_0_bits_control; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_CarryDepenIn_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_CarryDepenIn_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire [31:0] Loop_2_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopExit_0_ready; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopExit_0_valid; // @[bbgemm.scala 66:22]
  wire [9:0] Loop_2_io_loopExit_0_bits_taskID; // @[bbgemm.scala 66:22]
  wire  Loop_2_io_loopExit_0_bits_control; // @[bbgemm.scala 66:22]
  wire  Loop_3_clock; // @[bbgemm.scala 68:22]
  wire  Loop_3_reset; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_enable_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_enable_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_enable_bits_taskID; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_enable_bits_control; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_0_valid; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_1_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_1_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_InLiveIn_1_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_1_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_2_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_2_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_InLiveIn_2_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_2_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_3_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_InLiveIn_3_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_InLiveIn_3_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_3_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field3_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_OutLiveIn_field3_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_activate_loop_start_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_activate_loop_start_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_activate_loop_start_bits_control; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_activate_loop_back_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_activate_loop_back_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_activate_loop_back_bits_control; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopBack_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopBack_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_loopBack_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopBack_0_bits_control; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopFinish_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopFinish_0_valid; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopFinish_0_bits_control; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_CarryDepenIn_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_CarryDepenIn_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire [31:0] Loop_3_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopExit_0_ready; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopExit_0_valid; // @[bbgemm.scala 68:22]
  wire [9:0] Loop_3_io_loopExit_0_bits_taskID; // @[bbgemm.scala 68:22]
  wire  Loop_3_io_loopExit_0_bits_control; // @[bbgemm.scala 68:22]
  wire  Loop_4_clock; // @[bbgemm.scala 70:22]
  wire  Loop_4_reset; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_enable_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_enable_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_enable_bits_taskID; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_enable_bits_control; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_InLiveIn_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_InLiveIn_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_InLiveIn_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_0_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_InLiveIn_1_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_InLiveIn_1_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_InLiveIn_1_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_1_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_InLiveIn_2_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_InLiveIn_2_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_InLiveIn_2_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_2_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field2_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field1_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field0_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_OutLiveIn_field0_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_activate_loop_start_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_activate_loop_start_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_activate_loop_start_bits_control; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_activate_loop_back_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_activate_loop_back_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_activate_loop_back_bits_control; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopBack_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopBack_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_loopBack_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopBack_0_bits_control; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopFinish_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopFinish_0_valid; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopFinish_0_bits_control; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_CarryDepenIn_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_CarryDepenIn_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_CarryDepenIn_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_CarryDepenIn_0_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_CarryDepenOut_field0_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire [31:0] Loop_4_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopExit_0_ready; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopExit_0_valid; // @[bbgemm.scala 70:22]
  wire [9:0] Loop_4_io_loopExit_0_bits_taskID; // @[bbgemm.scala 70:22]
  wire  Loop_4_io_loopExit_0_bits_control; // @[bbgemm.scala 70:22]
  wire  bb_0_clock; // @[bbgemm.scala 78:20]
  wire  bb_0_reset; // @[bbgemm.scala 78:20]
  wire  bb_0_io_predicateIn_0_ready; // @[bbgemm.scala 78:20]
  wire  bb_0_io_predicateIn_0_valid; // @[bbgemm.scala 78:20]
  wire [9:0] bb_0_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 78:20]
  wire  bb_0_io_predicateIn_0_bits_control; // @[bbgemm.scala 78:20]
  wire  bb_0_io_Out_0_ready; // @[bbgemm.scala 78:20]
  wire  bb_0_io_Out_0_valid; // @[bbgemm.scala 78:20]
  wire [9:0] bb_0_io_Out_0_bits_taskID; // @[bbgemm.scala 78:20]
  wire  bb_0_io_Out_0_bits_control; // @[bbgemm.scala 78:20]
  wire  bb_1_clock; // @[bbgemm.scala 80:20]
  wire  bb_1_reset; // @[bbgemm.scala 80:20]
  wire  bb_1_io_MaskBB_0_ready; // @[bbgemm.scala 80:20]
  wire  bb_1_io_MaskBB_0_valid; // @[bbgemm.scala 80:20]
  wire [1:0] bb_1_io_MaskBB_0_bits; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_0_ready; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_0_valid; // @[bbgemm.scala 80:20]
  wire [9:0] bb_1_io_Out_0_bits_taskID; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_1_ready; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_1_valid; // @[bbgemm.scala 80:20]
  wire [9:0] bb_1_io_Out_1_bits_taskID; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_1_bits_control; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_2_ready; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_2_valid; // @[bbgemm.scala 80:20]
  wire [9:0] bb_1_io_Out_2_bits_taskID; // @[bbgemm.scala 80:20]
  wire  bb_1_io_Out_2_bits_control; // @[bbgemm.scala 80:20]
  wire  bb_1_io_predicateIn_0_ready; // @[bbgemm.scala 80:20]
  wire  bb_1_io_predicateIn_0_valid; // @[bbgemm.scala 80:20]
  wire [9:0] bb_1_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 80:20]
  wire  bb_1_io_predicateIn_0_bits_control; // @[bbgemm.scala 80:20]
  wire  bb_1_io_predicateIn_1_ready; // @[bbgemm.scala 80:20]
  wire  bb_1_io_predicateIn_1_valid; // @[bbgemm.scala 80:20]
  wire [9:0] bb_1_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 80:20]
  wire  bb_1_io_predicateIn_1_bits_control; // @[bbgemm.scala 80:20]
  wire  bb_2_clock; // @[bbgemm.scala 82:20]
  wire  bb_2_reset; // @[bbgemm.scala 82:20]
  wire  bb_2_io_MaskBB_0_ready; // @[bbgemm.scala 82:20]
  wire  bb_2_io_MaskBB_0_valid; // @[bbgemm.scala 82:20]
  wire [1:0] bb_2_io_MaskBB_0_bits; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_0_ready; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_0_valid; // @[bbgemm.scala 82:20]
  wire [9:0] bb_2_io_Out_0_bits_taskID; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_1_ready; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_1_valid; // @[bbgemm.scala 82:20]
  wire [9:0] bb_2_io_Out_1_bits_taskID; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_1_bits_control; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_2_ready; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_2_valid; // @[bbgemm.scala 82:20]
  wire [9:0] bb_2_io_Out_2_bits_taskID; // @[bbgemm.scala 82:20]
  wire  bb_2_io_Out_2_bits_control; // @[bbgemm.scala 82:20]
  wire  bb_2_io_predicateIn_0_ready; // @[bbgemm.scala 82:20]
  wire  bb_2_io_predicateIn_0_valid; // @[bbgemm.scala 82:20]
  wire [9:0] bb_2_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 82:20]
  wire  bb_2_io_predicateIn_0_bits_control; // @[bbgemm.scala 82:20]
  wire  bb_2_io_predicateIn_1_ready; // @[bbgemm.scala 82:20]
  wire  bb_2_io_predicateIn_1_valid; // @[bbgemm.scala 82:20]
  wire [9:0] bb_2_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 82:20]
  wire  bb_2_io_predicateIn_1_bits_control; // @[bbgemm.scala 82:20]
  wire  bb_3_clock; // @[bbgemm.scala 84:20]
  wire  bb_3_reset; // @[bbgemm.scala 84:20]
  wire  bb_3_io_MaskBB_0_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_MaskBB_0_valid; // @[bbgemm.scala 84:20]
  wire [1:0] bb_3_io_MaskBB_0_bits; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_0_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_0_valid; // @[bbgemm.scala 84:20]
  wire [9:0] bb_3_io_Out_0_bits_taskID; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_1_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_1_valid; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_2_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_2_valid; // @[bbgemm.scala 84:20]
  wire [9:0] bb_3_io_Out_2_bits_taskID; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_2_bits_control; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_3_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_3_valid; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_3_bits_control; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_4_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_4_valid; // @[bbgemm.scala 84:20]
  wire [9:0] bb_3_io_Out_4_bits_taskID; // @[bbgemm.scala 84:20]
  wire  bb_3_io_Out_4_bits_control; // @[bbgemm.scala 84:20]
  wire  bb_3_io_predicateIn_0_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_predicateIn_0_valid; // @[bbgemm.scala 84:20]
  wire [9:0] bb_3_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 84:20]
  wire  bb_3_io_predicateIn_0_bits_control; // @[bbgemm.scala 84:20]
  wire  bb_3_io_predicateIn_1_ready; // @[bbgemm.scala 84:20]
  wire  bb_3_io_predicateIn_1_valid; // @[bbgemm.scala 84:20]
  wire [9:0] bb_3_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 84:20]
  wire  bb_3_io_predicateIn_1_bits_control; // @[bbgemm.scala 84:20]
  wire  bb_4_clock; // @[bbgemm.scala 86:20]
  wire  bb_4_reset; // @[bbgemm.scala 86:20]
  wire  bb_4_io_MaskBB_0_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_MaskBB_0_valid; // @[bbgemm.scala 86:20]
  wire [1:0] bb_4_io_MaskBB_0_bits; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_0_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_0_valid; // @[bbgemm.scala 86:20]
  wire [9:0] bb_4_io_Out_0_bits_taskID; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_1_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_1_valid; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_2_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_2_valid; // @[bbgemm.scala 86:20]
  wire [9:0] bb_4_io_Out_2_bits_taskID; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_2_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_3_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_3_valid; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_3_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_4_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_4_valid; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_4_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_5_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_5_valid; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_5_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_6_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_6_valid; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_6_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_7_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_7_valid; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_7_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_8_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_8_valid; // @[bbgemm.scala 86:20]
  wire [9:0] bb_4_io_Out_8_bits_taskID; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_8_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_9_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_9_valid; // @[bbgemm.scala 86:20]
  wire [9:0] bb_4_io_Out_9_bits_taskID; // @[bbgemm.scala 86:20]
  wire  bb_4_io_Out_9_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_predicateIn_0_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_predicateIn_0_valid; // @[bbgemm.scala 86:20]
  wire [9:0] bb_4_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 86:20]
  wire  bb_4_io_predicateIn_0_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_4_io_predicateIn_1_ready; // @[bbgemm.scala 86:20]
  wire  bb_4_io_predicateIn_1_valid; // @[bbgemm.scala 86:20]
  wire [9:0] bb_4_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 86:20]
  wire  bb_4_io_predicateIn_1_bits_control; // @[bbgemm.scala 86:20]
  wire  bb_5_clock; // @[bbgemm.scala 88:20]
  wire  bb_5_reset; // @[bbgemm.scala 88:20]
  wire  bb_5_io_MaskBB_0_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_MaskBB_0_valid; // @[bbgemm.scala 88:20]
  wire [1:0] bb_5_io_MaskBB_0_bits; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_0_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_0_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_0_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_1_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_1_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_1_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_2_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_2_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_2_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_3_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_3_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_3_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_3_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_4_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_4_valid; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_4_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_5_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_5_valid; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_5_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_6_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_6_valid; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_6_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_7_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_7_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_7_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_7_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_8_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_8_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_8_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_8_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_9_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_9_valid; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_9_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_10_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_10_valid; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_10_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_11_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_11_valid; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_11_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_12_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_12_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_12_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_12_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_13_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_13_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_13_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_13_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_14_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_14_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_14_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_14_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_15_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_15_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_15_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_15_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_16_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_16_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_16_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_16_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_17_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_17_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_Out_17_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_Out_17_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_predicateIn_0_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_predicateIn_0_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_predicateIn_0_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_5_io_predicateIn_1_ready; // @[bbgemm.scala 88:20]
  wire  bb_5_io_predicateIn_1_valid; // @[bbgemm.scala 88:20]
  wire [9:0] bb_5_io_predicateIn_1_bits_taskID; // @[bbgemm.scala 88:20]
  wire  bb_5_io_predicateIn_1_bits_control; // @[bbgemm.scala 88:20]
  wire  bb_6_clock; // @[bbgemm.scala 90:20]
  wire  bb_6_reset; // @[bbgemm.scala 90:20]
  wire  bb_6_io_predicateIn_0_ready; // @[bbgemm.scala 90:20]
  wire  bb_6_io_predicateIn_0_valid; // @[bbgemm.scala 90:20]
  wire [9:0] bb_6_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 90:20]
  wire  bb_6_io_predicateIn_0_bits_control; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_0_ready; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_0_valid; // @[bbgemm.scala 90:20]
  wire [9:0] bb_6_io_Out_0_bits_taskID; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_1_ready; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_1_valid; // @[bbgemm.scala 90:20]
  wire [9:0] bb_6_io_Out_1_bits_taskID; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_2_ready; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_2_valid; // @[bbgemm.scala 90:20]
  wire [9:0] bb_6_io_Out_2_bits_taskID; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_2_bits_control; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_3_ready; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_3_valid; // @[bbgemm.scala 90:20]
  wire [9:0] bb_6_io_Out_3_bits_taskID; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_3_bits_control; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_4_ready; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_4_valid; // @[bbgemm.scala 90:20]
  wire [9:0] bb_6_io_Out_4_bits_taskID; // @[bbgemm.scala 90:20]
  wire  bb_6_io_Out_4_bits_control; // @[bbgemm.scala 90:20]
  wire  bb_7_clock; // @[bbgemm.scala 92:20]
  wire  bb_7_reset; // @[bbgemm.scala 92:20]
  wire  bb_7_io_predicateIn_0_ready; // @[bbgemm.scala 92:20]
  wire  bb_7_io_predicateIn_0_valid; // @[bbgemm.scala 92:20]
  wire [9:0] bb_7_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 92:20]
  wire  bb_7_io_predicateIn_0_bits_control; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_0_ready; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_0_valid; // @[bbgemm.scala 92:20]
  wire [9:0] bb_7_io_Out_0_bits_taskID; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_1_ready; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_1_valid; // @[bbgemm.scala 92:20]
  wire [9:0] bb_7_io_Out_1_bits_taskID; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_2_ready; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_2_valid; // @[bbgemm.scala 92:20]
  wire [9:0] bb_7_io_Out_2_bits_taskID; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_2_bits_control; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_3_ready; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_3_valid; // @[bbgemm.scala 92:20]
  wire [9:0] bb_7_io_Out_3_bits_taskID; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_3_bits_control; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_4_ready; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_4_valid; // @[bbgemm.scala 92:20]
  wire [9:0] bb_7_io_Out_4_bits_taskID; // @[bbgemm.scala 92:20]
  wire  bb_7_io_Out_4_bits_control; // @[bbgemm.scala 92:20]
  wire  bb_8_clock; // @[bbgemm.scala 94:20]
  wire  bb_8_reset; // @[bbgemm.scala 94:20]
  wire  bb_8_io_predicateIn_0_ready; // @[bbgemm.scala 94:20]
  wire  bb_8_io_predicateIn_0_valid; // @[bbgemm.scala 94:20]
  wire [9:0] bb_8_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 94:20]
  wire  bb_8_io_predicateIn_0_bits_control; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_0_ready; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_0_valid; // @[bbgemm.scala 94:20]
  wire [9:0] bb_8_io_Out_0_bits_taskID; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_1_ready; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_1_valid; // @[bbgemm.scala 94:20]
  wire [9:0] bb_8_io_Out_1_bits_taskID; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_2_ready; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_2_valid; // @[bbgemm.scala 94:20]
  wire [9:0] bb_8_io_Out_2_bits_taskID; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_2_bits_control; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_3_ready; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_3_valid; // @[bbgemm.scala 94:20]
  wire [9:0] bb_8_io_Out_3_bits_taskID; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_3_bits_control; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_4_ready; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_4_valid; // @[bbgemm.scala 94:20]
  wire [9:0] bb_8_io_Out_4_bits_taskID; // @[bbgemm.scala 94:20]
  wire  bb_8_io_Out_4_bits_control; // @[bbgemm.scala 94:20]
  wire  bb_9_clock; // @[bbgemm.scala 96:20]
  wire  bb_9_reset; // @[bbgemm.scala 96:20]
  wire  bb_9_io_predicateIn_0_ready; // @[bbgemm.scala 96:20]
  wire  bb_9_io_predicateIn_0_valid; // @[bbgemm.scala 96:20]
  wire [9:0] bb_9_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 96:20]
  wire  bb_9_io_predicateIn_0_bits_control; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_0_ready; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_0_valid; // @[bbgemm.scala 96:20]
  wire [9:0] bb_9_io_Out_0_bits_taskID; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_1_ready; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_1_valid; // @[bbgemm.scala 96:20]
  wire [9:0] bb_9_io_Out_1_bits_taskID; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_2_ready; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_2_valid; // @[bbgemm.scala 96:20]
  wire [9:0] bb_9_io_Out_2_bits_taskID; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_2_bits_control; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_3_ready; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_3_valid; // @[bbgemm.scala 96:20]
  wire [9:0] bb_9_io_Out_3_bits_taskID; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_3_bits_control; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_4_ready; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_4_valid; // @[bbgemm.scala 96:20]
  wire [9:0] bb_9_io_Out_4_bits_taskID; // @[bbgemm.scala 96:20]
  wire  bb_9_io_Out_4_bits_control; // @[bbgemm.scala 96:20]
  wire  bb_10_clock; // @[bbgemm.scala 98:21]
  wire  bb_10_reset; // @[bbgemm.scala 98:21]
  wire  bb_10_io_predicateIn_0_ready; // @[bbgemm.scala 98:21]
  wire  bb_10_io_predicateIn_0_valid; // @[bbgemm.scala 98:21]
  wire [9:0] bb_10_io_predicateIn_0_bits_taskID; // @[bbgemm.scala 98:21]
  wire  bb_10_io_predicateIn_0_bits_control; // @[bbgemm.scala 98:21]
  wire  bb_10_io_Out_0_ready; // @[bbgemm.scala 98:21]
  wire  bb_10_io_Out_0_valid; // @[bbgemm.scala 98:21]
  wire [9:0] bb_10_io_Out_0_bits_taskID; // @[bbgemm.scala 98:21]
  wire  bb_10_io_Out_0_bits_control; // @[bbgemm.scala 98:21]
  wire  br_0_clock; // @[bbgemm.scala 107:20]
  wire  br_0_reset; // @[bbgemm.scala 107:20]
  wire  br_0_io_enable_ready; // @[bbgemm.scala 107:20]
  wire  br_0_io_enable_valid; // @[bbgemm.scala 107:20]
  wire [9:0] br_0_io_enable_bits_taskID; // @[bbgemm.scala 107:20]
  wire  br_0_io_enable_bits_control; // @[bbgemm.scala 107:20]
  wire  br_0_io_Out_0_ready; // @[bbgemm.scala 107:20]
  wire  br_0_io_Out_0_valid; // @[bbgemm.scala 107:20]
  wire [9:0] br_0_io_Out_0_bits_taskID; // @[bbgemm.scala 107:20]
  wire  br_0_io_Out_0_bits_control; // @[bbgemm.scala 107:20]
  wire  phi1_clock; // @[bbgemm.scala 110:20]
  wire  phi1_reset; // @[bbgemm.scala 110:20]
  wire  phi1_io_enable_ready; // @[bbgemm.scala 110:20]
  wire  phi1_io_enable_valid; // @[bbgemm.scala 110:20]
  wire [9:0] phi1_io_enable_bits_taskID; // @[bbgemm.scala 110:20]
  wire  phi1_io_enable_bits_control; // @[bbgemm.scala 110:20]
  wire  phi1_io_InData_0_ready; // @[bbgemm.scala 110:20]
  wire  phi1_io_InData_0_valid; // @[bbgemm.scala 110:20]
  wire [9:0] phi1_io_InData_0_bits_taskID; // @[bbgemm.scala 110:20]
  wire  phi1_io_InData_1_ready; // @[bbgemm.scala 110:20]
  wire  phi1_io_InData_1_valid; // @[bbgemm.scala 110:20]
  wire [9:0] phi1_io_InData_1_bits_taskID; // @[bbgemm.scala 110:20]
  wire [31:0] phi1_io_InData_1_bits_data; // @[bbgemm.scala 110:20]
  wire  phi1_io_Mask_ready; // @[bbgemm.scala 110:20]
  wire  phi1_io_Mask_valid; // @[bbgemm.scala 110:20]
  wire [1:0] phi1_io_Mask_bits; // @[bbgemm.scala 110:20]
  wire  phi1_io_Out_0_ready; // @[bbgemm.scala 110:20]
  wire  phi1_io_Out_0_valid; // @[bbgemm.scala 110:20]
  wire [31:0] phi1_io_Out_0_bits_data; // @[bbgemm.scala 110:20]
  wire  phi1_io_Out_1_ready; // @[bbgemm.scala 110:20]
  wire  phi1_io_Out_1_valid; // @[bbgemm.scala 110:20]
  wire [9:0] phi1_io_Out_1_bits_taskID; // @[bbgemm.scala 110:20]
  wire [31:0] phi1_io_Out_1_bits_data; // @[bbgemm.scala 110:20]
  wire  br_2_clock; // @[bbgemm.scala 113:20]
  wire  br_2_reset; // @[bbgemm.scala 113:20]
  wire  br_2_io_enable_ready; // @[bbgemm.scala 113:20]
  wire  br_2_io_enable_valid; // @[bbgemm.scala 113:20]
  wire [9:0] br_2_io_enable_bits_taskID; // @[bbgemm.scala 113:20]
  wire  br_2_io_enable_bits_control; // @[bbgemm.scala 113:20]
  wire  br_2_io_Out_0_ready; // @[bbgemm.scala 113:20]
  wire  br_2_io_Out_0_valid; // @[bbgemm.scala 113:20]
  wire [9:0] br_2_io_Out_0_bits_taskID; // @[bbgemm.scala 113:20]
  wire  br_2_io_Out_0_bits_control; // @[bbgemm.scala 113:20]
  wire  phi3_clock; // @[bbgemm.scala 116:20]
  wire  phi3_reset; // @[bbgemm.scala 116:20]
  wire  phi3_io_enable_ready; // @[bbgemm.scala 116:20]
  wire  phi3_io_enable_valid; // @[bbgemm.scala 116:20]
  wire [9:0] phi3_io_enable_bits_taskID; // @[bbgemm.scala 116:20]
  wire  phi3_io_enable_bits_control; // @[bbgemm.scala 116:20]
  wire  phi3_io_InData_0_ready; // @[bbgemm.scala 116:20]
  wire  phi3_io_InData_0_valid; // @[bbgemm.scala 116:20]
  wire [9:0] phi3_io_InData_0_bits_taskID; // @[bbgemm.scala 116:20]
  wire  phi3_io_InData_1_ready; // @[bbgemm.scala 116:20]
  wire  phi3_io_InData_1_valid; // @[bbgemm.scala 116:20]
  wire [9:0] phi3_io_InData_1_bits_taskID; // @[bbgemm.scala 116:20]
  wire [31:0] phi3_io_InData_1_bits_data; // @[bbgemm.scala 116:20]
  wire  phi3_io_Mask_ready; // @[bbgemm.scala 116:20]
  wire  phi3_io_Mask_valid; // @[bbgemm.scala 116:20]
  wire [1:0] phi3_io_Mask_bits; // @[bbgemm.scala 116:20]
  wire  phi3_io_Out_0_ready; // @[bbgemm.scala 116:20]
  wire  phi3_io_Out_0_valid; // @[bbgemm.scala 116:20]
  wire [31:0] phi3_io_Out_0_bits_data; // @[bbgemm.scala 116:20]
  wire  phi3_io_Out_1_ready; // @[bbgemm.scala 116:20]
  wire  phi3_io_Out_1_valid; // @[bbgemm.scala 116:20]
  wire [9:0] phi3_io_Out_1_bits_taskID; // @[bbgemm.scala 116:20]
  wire [31:0] phi3_io_Out_1_bits_data; // @[bbgemm.scala 116:20]
  wire  br_4_clock; // @[bbgemm.scala 119:20]
  wire  br_4_reset; // @[bbgemm.scala 119:20]
  wire  br_4_io_enable_ready; // @[bbgemm.scala 119:20]
  wire  br_4_io_enable_valid; // @[bbgemm.scala 119:20]
  wire [9:0] br_4_io_enable_bits_taskID; // @[bbgemm.scala 119:20]
  wire  br_4_io_enable_bits_control; // @[bbgemm.scala 119:20]
  wire  br_4_io_Out_0_ready; // @[bbgemm.scala 119:20]
  wire  br_4_io_Out_0_valid; // @[bbgemm.scala 119:20]
  wire [9:0] br_4_io_Out_0_bits_taskID; // @[bbgemm.scala 119:20]
  wire  br_4_io_Out_0_bits_control; // @[bbgemm.scala 119:20]
  wire  phi5_clock; // @[bbgemm.scala 122:20]
  wire  phi5_reset; // @[bbgemm.scala 122:20]
  wire  phi5_io_enable_ready; // @[bbgemm.scala 122:20]
  wire  phi5_io_enable_valid; // @[bbgemm.scala 122:20]
  wire [9:0] phi5_io_enable_bits_taskID; // @[bbgemm.scala 122:20]
  wire  phi5_io_enable_bits_control; // @[bbgemm.scala 122:20]
  wire  phi5_io_InData_0_ready; // @[bbgemm.scala 122:20]
  wire  phi5_io_InData_0_valid; // @[bbgemm.scala 122:20]
  wire [9:0] phi5_io_InData_0_bits_taskID; // @[bbgemm.scala 122:20]
  wire  phi5_io_InData_1_ready; // @[bbgemm.scala 122:20]
  wire  phi5_io_InData_1_valid; // @[bbgemm.scala 122:20]
  wire [9:0] phi5_io_InData_1_bits_taskID; // @[bbgemm.scala 122:20]
  wire [31:0] phi5_io_InData_1_bits_data; // @[bbgemm.scala 122:20]
  wire  phi5_io_Mask_ready; // @[bbgemm.scala 122:20]
  wire  phi5_io_Mask_valid; // @[bbgemm.scala 122:20]
  wire [1:0] phi5_io_Mask_bits; // @[bbgemm.scala 122:20]
  wire  phi5_io_Out_0_ready; // @[bbgemm.scala 122:20]
  wire  phi5_io_Out_0_valid; // @[bbgemm.scala 122:20]
  wire [31:0] phi5_io_Out_0_bits_data; // @[bbgemm.scala 122:20]
  wire  phi5_io_Out_1_ready; // @[bbgemm.scala 122:20]
  wire  phi5_io_Out_1_valid; // @[bbgemm.scala 122:20]
  wire [9:0] phi5_io_Out_1_bits_taskID; // @[bbgemm.scala 122:20]
  wire [31:0] phi5_io_Out_1_bits_data; // @[bbgemm.scala 122:20]
  wire  binaryOp_6_clock; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_reset; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_enable_ready; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_enable_valid; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_enable_bits_control; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_Out_0_ready; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_Out_0_valid; // @[bbgemm.scala 125:26]
  wire [31:0] binaryOp_6_io_Out_0_bits_data; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_LeftIO_ready; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_LeftIO_valid; // @[bbgemm.scala 125:26]
  wire [31:0] binaryOp_6_io_LeftIO_bits_data; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_RightIO_ready; // @[bbgemm.scala 125:26]
  wire  binaryOp_6_io_RightIO_valid; // @[bbgemm.scala 125:26]
  wire  br_7_clock; // @[bbgemm.scala 128:20]
  wire  br_7_reset; // @[bbgemm.scala 128:20]
  wire  br_7_io_enable_ready; // @[bbgemm.scala 128:20]
  wire  br_7_io_enable_valid; // @[bbgemm.scala 128:20]
  wire [9:0] br_7_io_enable_bits_taskID; // @[bbgemm.scala 128:20]
  wire  br_7_io_enable_bits_control; // @[bbgemm.scala 128:20]
  wire  br_7_io_Out_0_ready; // @[bbgemm.scala 128:20]
  wire  br_7_io_Out_0_valid; // @[bbgemm.scala 128:20]
  wire [9:0] br_7_io_Out_0_bits_taskID; // @[bbgemm.scala 128:20]
  wire  br_7_io_Out_0_bits_control; // @[bbgemm.scala 128:20]
  wire  phi8_clock; // @[bbgemm.scala 131:20]
  wire  phi8_reset; // @[bbgemm.scala 131:20]
  wire  phi8_io_enable_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_enable_valid; // @[bbgemm.scala 131:20]
  wire [9:0] phi8_io_enable_bits_taskID; // @[bbgemm.scala 131:20]
  wire  phi8_io_enable_bits_control; // @[bbgemm.scala 131:20]
  wire  phi8_io_InData_0_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_InData_0_valid; // @[bbgemm.scala 131:20]
  wire [9:0] phi8_io_InData_0_bits_taskID; // @[bbgemm.scala 131:20]
  wire  phi8_io_InData_1_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_InData_1_valid; // @[bbgemm.scala 131:20]
  wire [9:0] phi8_io_InData_1_bits_taskID; // @[bbgemm.scala 131:20]
  wire [31:0] phi8_io_InData_1_bits_data; // @[bbgemm.scala 131:20]
  wire  phi8_io_Mask_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_Mask_valid; // @[bbgemm.scala 131:20]
  wire [1:0] phi8_io_Mask_bits; // @[bbgemm.scala 131:20]
  wire  phi8_io_Out_0_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_Out_0_valid; // @[bbgemm.scala 131:20]
  wire [31:0] phi8_io_Out_0_bits_data; // @[bbgemm.scala 131:20]
  wire  phi8_io_Out_1_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_Out_1_valid; // @[bbgemm.scala 131:20]
  wire [31:0] phi8_io_Out_1_bits_data; // @[bbgemm.scala 131:20]
  wire  phi8_io_Out_2_ready; // @[bbgemm.scala 131:20]
  wire  phi8_io_Out_2_valid; // @[bbgemm.scala 131:20]
  wire [9:0] phi8_io_Out_2_bits_taskID; // @[bbgemm.scala 131:20]
  wire [31:0] phi8_io_Out_2_bits_data; // @[bbgemm.scala 131:20]
  wire  binaryOp_9_clock; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_reset; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_enable_ready; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_enable_valid; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_enable_bits_control; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_Out_0_ready; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_Out_0_valid; // @[bbgemm.scala 134:26]
  wire [31:0] binaryOp_9_io_Out_0_bits_data; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_LeftIO_ready; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_LeftIO_valid; // @[bbgemm.scala 134:26]
  wire [31:0] binaryOp_9_io_LeftIO_bits_data; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_RightIO_ready; // @[bbgemm.scala 134:26]
  wire  binaryOp_9_io_RightIO_valid; // @[bbgemm.scala 134:26]
  wire [31:0] binaryOp_9_io_RightIO_bits_data; // @[bbgemm.scala 134:26]
  wire  binaryOp_10_clock; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_reset; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_enable_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_enable_valid; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_enable_bits_control; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_Out_0_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_Out_0_valid; // @[bbgemm.scala 137:27]
  wire [31:0] binaryOp_10_io_Out_0_bits_data; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_LeftIO_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_LeftIO_valid; // @[bbgemm.scala 137:27]
  wire [31:0] binaryOp_10_io_LeftIO_bits_data; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_RightIO_ready; // @[bbgemm.scala 137:27]
  wire  binaryOp_10_io_RightIO_valid; // @[bbgemm.scala 137:27]
  wire  binaryOp_11_clock; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_reset; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_enable_ready; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_enable_valid; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_enable_bits_control; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_Out_0_ready; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_Out_0_valid; // @[bbgemm.scala 140:27]
  wire [31:0] binaryOp_11_io_Out_0_bits_data; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_LeftIO_ready; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_LeftIO_valid; // @[bbgemm.scala 140:27]
  wire [31:0] binaryOp_11_io_LeftIO_bits_data; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_RightIO_ready; // @[bbgemm.scala 140:27]
  wire  binaryOp_11_io_RightIO_valid; // @[bbgemm.scala 140:27]
  wire [31:0] binaryOp_11_io_RightIO_bits_data; // @[bbgemm.scala 140:27]
  wire  binaryOp_12_clock; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_reset; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_enable_ready; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_enable_valid; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_enable_bits_control; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_Out_0_ready; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_Out_0_valid; // @[bbgemm.scala 143:27]
  wire [31:0] binaryOp_12_io_Out_0_bits_data; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_LeftIO_ready; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_LeftIO_valid; // @[bbgemm.scala 143:27]
  wire [31:0] binaryOp_12_io_LeftIO_bits_data; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_RightIO_ready; // @[bbgemm.scala 143:27]
  wire  binaryOp_12_io_RightIO_valid; // @[bbgemm.scala 143:27]
  wire [31:0] binaryOp_12_io_RightIO_bits_data; // @[bbgemm.scala 143:27]
  wire  Gep_13_clock; // @[bbgemm.scala 146:22]
  wire  Gep_13_reset; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_enable_ready; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_enable_valid; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_enable_bits_control; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_Out_0_ready; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_Out_0_valid; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_Out_0_bits_predicate; // @[bbgemm.scala 146:22]
  wire [9:0] Gep_13_io_Out_0_bits_taskID; // @[bbgemm.scala 146:22]
  wire [31:0] Gep_13_io_Out_0_bits_data; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_baseAddress_ready; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_baseAddress_valid; // @[bbgemm.scala 146:22]
  wire [9:0] Gep_13_io_baseAddress_bits_taskID; // @[bbgemm.scala 146:22]
  wire [31:0] Gep_13_io_baseAddress_bits_data; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_idx_0_ready; // @[bbgemm.scala 146:22]
  wire  Gep_13_io_idx_0_valid; // @[bbgemm.scala 146:22]
  wire [31:0] Gep_13_io_idx_0_bits_data; // @[bbgemm.scala 146:22]
  wire  ld_14_clock; // @[bbgemm.scala 149:21]
  wire  ld_14_reset; // @[bbgemm.scala 149:21]
  wire  ld_14_io_enable_ready; // @[bbgemm.scala 149:21]
  wire  ld_14_io_enable_valid; // @[bbgemm.scala 149:21]
  wire [9:0] ld_14_io_enable_bits_taskID; // @[bbgemm.scala 149:21]
  wire  ld_14_io_enable_bits_control; // @[bbgemm.scala 149:21]
  wire  ld_14_io_Out_0_ready; // @[bbgemm.scala 149:21]
  wire  ld_14_io_Out_0_valid; // @[bbgemm.scala 149:21]
  wire [9:0] ld_14_io_Out_0_bits_taskID; // @[bbgemm.scala 149:21]
  wire [31:0] ld_14_io_Out_0_bits_data; // @[bbgemm.scala 149:21]
  wire  ld_14_io_GepAddr_ready; // @[bbgemm.scala 149:21]
  wire  ld_14_io_GepAddr_valid; // @[bbgemm.scala 149:21]
  wire  ld_14_io_GepAddr_bits_predicate; // @[bbgemm.scala 149:21]
  wire [9:0] ld_14_io_GepAddr_bits_taskID; // @[bbgemm.scala 149:21]
  wire [31:0] ld_14_io_GepAddr_bits_data; // @[bbgemm.scala 149:21]
  wire  ld_14_io_memReq_ready; // @[bbgemm.scala 149:21]
  wire  ld_14_io_memReq_valid; // @[bbgemm.scala 149:21]
  wire [31:0] ld_14_io_memReq_bits_address; // @[bbgemm.scala 149:21]
  wire [9:0] ld_14_io_memReq_bits_taskID; // @[bbgemm.scala 149:21]
  wire  ld_14_io_memResp_valid; // @[bbgemm.scala 149:21]
  wire [31:0] ld_14_io_memResp_data; // @[bbgemm.scala 149:21]
  wire  br_15_clock; // @[bbgemm.scala 152:21]
  wire  br_15_reset; // @[bbgemm.scala 152:21]
  wire  br_15_io_enable_ready; // @[bbgemm.scala 152:21]
  wire  br_15_io_enable_valid; // @[bbgemm.scala 152:21]
  wire [9:0] br_15_io_enable_bits_taskID; // @[bbgemm.scala 152:21]
  wire  br_15_io_enable_bits_control; // @[bbgemm.scala 152:21]
  wire  br_15_io_Out_0_ready; // @[bbgemm.scala 152:21]
  wire  br_15_io_Out_0_valid; // @[bbgemm.scala 152:21]
  wire [9:0] br_15_io_Out_0_bits_taskID; // @[bbgemm.scala 152:21]
  wire  br_15_io_Out_0_bits_control; // @[bbgemm.scala 152:21]
  wire  phi16_clock; // @[bbgemm.scala 155:21]
  wire  phi16_reset; // @[bbgemm.scala 155:21]
  wire  phi16_io_enable_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_enable_valid; // @[bbgemm.scala 155:21]
  wire [9:0] phi16_io_enable_bits_taskID; // @[bbgemm.scala 155:21]
  wire  phi16_io_enable_bits_control; // @[bbgemm.scala 155:21]
  wire  phi16_io_InData_0_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_InData_0_valid; // @[bbgemm.scala 155:21]
  wire [9:0] phi16_io_InData_0_bits_taskID; // @[bbgemm.scala 155:21]
  wire  phi16_io_InData_1_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_InData_1_valid; // @[bbgemm.scala 155:21]
  wire [9:0] phi16_io_InData_1_bits_taskID; // @[bbgemm.scala 155:21]
  wire [31:0] phi16_io_InData_1_bits_data; // @[bbgemm.scala 155:21]
  wire  phi16_io_Mask_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_Mask_valid; // @[bbgemm.scala 155:21]
  wire [1:0] phi16_io_Mask_bits; // @[bbgemm.scala 155:21]
  wire  phi16_io_Out_0_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_Out_0_valid; // @[bbgemm.scala 155:21]
  wire [31:0] phi16_io_Out_0_bits_data; // @[bbgemm.scala 155:21]
  wire  phi16_io_Out_1_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_Out_1_valid; // @[bbgemm.scala 155:21]
  wire [31:0] phi16_io_Out_1_bits_data; // @[bbgemm.scala 155:21]
  wire  phi16_io_Out_2_ready; // @[bbgemm.scala 155:21]
  wire  phi16_io_Out_2_valid; // @[bbgemm.scala 155:21]
  wire [9:0] phi16_io_Out_2_bits_taskID; // @[bbgemm.scala 155:21]
  wire [31:0] phi16_io_Out_2_bits_data; // @[bbgemm.scala 155:21]
  wire  binaryOp_17_clock; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_reset; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_enable_ready; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_enable_valid; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_enable_bits_control; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_Out_0_ready; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_Out_0_valid; // @[bbgemm.scala 158:27]
  wire [31:0] binaryOp_17_io_Out_0_bits_data; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_LeftIO_ready; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_LeftIO_valid; // @[bbgemm.scala 158:27]
  wire [31:0] binaryOp_17_io_LeftIO_bits_data; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_RightIO_ready; // @[bbgemm.scala 158:27]
  wire  binaryOp_17_io_RightIO_valid; // @[bbgemm.scala 158:27]
  wire [31:0] binaryOp_17_io_RightIO_bits_data; // @[bbgemm.scala 158:27]
  wire  binaryOp_18_clock; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_reset; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_enable_ready; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_enable_valid; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_enable_bits_control; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_Out_0_ready; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_Out_0_valid; // @[bbgemm.scala 161:27]
  wire [31:0] binaryOp_18_io_Out_0_bits_data; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_LeftIO_ready; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_LeftIO_valid; // @[bbgemm.scala 161:27]
  wire [31:0] binaryOp_18_io_LeftIO_bits_data; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_RightIO_ready; // @[bbgemm.scala 161:27]
  wire  binaryOp_18_io_RightIO_valid; // @[bbgemm.scala 161:27]
  wire [31:0] binaryOp_18_io_RightIO_bits_data; // @[bbgemm.scala 161:27]
  wire  Gep_19_clock; // @[bbgemm.scala 164:22]
  wire  Gep_19_reset; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_enable_ready; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_enable_valid; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_enable_bits_control; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_Out_0_ready; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_Out_0_valid; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_Out_0_bits_predicate; // @[bbgemm.scala 164:22]
  wire [9:0] Gep_19_io_Out_0_bits_taskID; // @[bbgemm.scala 164:22]
  wire [31:0] Gep_19_io_Out_0_bits_data; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_baseAddress_ready; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_baseAddress_valid; // @[bbgemm.scala 164:22]
  wire [9:0] Gep_19_io_baseAddress_bits_taskID; // @[bbgemm.scala 164:22]
  wire [31:0] Gep_19_io_baseAddress_bits_data; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_idx_0_ready; // @[bbgemm.scala 164:22]
  wire  Gep_19_io_idx_0_valid; // @[bbgemm.scala 164:22]
  wire [31:0] Gep_19_io_idx_0_bits_data; // @[bbgemm.scala 164:22]
  wire  ld_20_clock; // @[bbgemm.scala 167:21]
  wire  ld_20_reset; // @[bbgemm.scala 167:21]
  wire  ld_20_io_enable_ready; // @[bbgemm.scala 167:21]
  wire  ld_20_io_enable_valid; // @[bbgemm.scala 167:21]
  wire [9:0] ld_20_io_enable_bits_taskID; // @[bbgemm.scala 167:21]
  wire  ld_20_io_enable_bits_control; // @[bbgemm.scala 167:21]
  wire  ld_20_io_Out_0_ready; // @[bbgemm.scala 167:21]
  wire  ld_20_io_Out_0_valid; // @[bbgemm.scala 167:21]
  wire [9:0] ld_20_io_Out_0_bits_taskID; // @[bbgemm.scala 167:21]
  wire [31:0] ld_20_io_Out_0_bits_data; // @[bbgemm.scala 167:21]
  wire  ld_20_io_GepAddr_ready; // @[bbgemm.scala 167:21]
  wire  ld_20_io_GepAddr_valid; // @[bbgemm.scala 167:21]
  wire  ld_20_io_GepAddr_bits_predicate; // @[bbgemm.scala 167:21]
  wire [9:0] ld_20_io_GepAddr_bits_taskID; // @[bbgemm.scala 167:21]
  wire [31:0] ld_20_io_GepAddr_bits_data; // @[bbgemm.scala 167:21]
  wire  ld_20_io_memReq_ready; // @[bbgemm.scala 167:21]
  wire  ld_20_io_memReq_valid; // @[bbgemm.scala 167:21]
  wire [31:0] ld_20_io_memReq_bits_address; // @[bbgemm.scala 167:21]
  wire [9:0] ld_20_io_memReq_bits_taskID; // @[bbgemm.scala 167:21]
  wire  ld_20_io_memResp_valid; // @[bbgemm.scala 167:21]
  wire [31:0] ld_20_io_memResp_data; // @[bbgemm.scala 167:21]
  wire  FP_21_clock; // @[bbgemm.scala 171:21]
  wire  FP_21_reset; // @[bbgemm.scala 171:21]
  wire  FP_21_io_enable_ready; // @[bbgemm.scala 171:21]
  wire  FP_21_io_enable_valid; // @[bbgemm.scala 171:21]
  wire [9:0] FP_21_io_enable_bits_taskID; // @[bbgemm.scala 171:21]
  wire  FP_21_io_enable_bits_control; // @[bbgemm.scala 171:21]
  wire  FP_21_io_Out_0_ready; // @[bbgemm.scala 171:21]
  wire  FP_21_io_Out_0_valid; // @[bbgemm.scala 171:21]
  wire [9:0] FP_21_io_Out_0_bits_taskID; // @[bbgemm.scala 171:21]
  wire [31:0] FP_21_io_Out_0_bits_data; // @[bbgemm.scala 171:21]
  wire  FP_21_io_LeftIO_ready; // @[bbgemm.scala 171:21]
  wire  FP_21_io_LeftIO_valid; // @[bbgemm.scala 171:21]
  wire [9:0] FP_21_io_LeftIO_bits_taskID; // @[bbgemm.scala 171:21]
  wire [31:0] FP_21_io_LeftIO_bits_data; // @[bbgemm.scala 171:21]
  wire  FP_21_io_RightIO_ready; // @[bbgemm.scala 171:21]
  wire  FP_21_io_RightIO_valid; // @[bbgemm.scala 171:21]
  wire [9:0] FP_21_io_RightIO_bits_taskID; // @[bbgemm.scala 171:21]
  wire [31:0] FP_21_io_RightIO_bits_data; // @[bbgemm.scala 171:21]
  wire  binaryOp_22_clock; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_reset; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_enable_ready; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_enable_valid; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_enable_bits_control; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_Out_0_ready; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_Out_0_valid; // @[bbgemm.scala 174:27]
  wire [31:0] binaryOp_22_io_Out_0_bits_data; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_LeftIO_ready; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_LeftIO_valid; // @[bbgemm.scala 174:27]
  wire [31:0] binaryOp_22_io_LeftIO_bits_data; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_RightIO_ready; // @[bbgemm.scala 174:27]
  wire  binaryOp_22_io_RightIO_valid; // @[bbgemm.scala 174:27]
  wire [31:0] binaryOp_22_io_RightIO_bits_data; // @[bbgemm.scala 174:27]
  wire  binaryOp_23_clock; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_reset; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_enable_ready; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_enable_valid; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_enable_bits_control; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_Out_0_ready; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_Out_0_valid; // @[bbgemm.scala 177:27]
  wire [31:0] binaryOp_23_io_Out_0_bits_data; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_LeftIO_ready; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_LeftIO_valid; // @[bbgemm.scala 177:27]
  wire [31:0] binaryOp_23_io_LeftIO_bits_data; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_RightIO_ready; // @[bbgemm.scala 177:27]
  wire  binaryOp_23_io_RightIO_valid; // @[bbgemm.scala 177:27]
  wire [31:0] binaryOp_23_io_RightIO_bits_data; // @[bbgemm.scala 177:27]
  wire  Gep_24_clock; // @[bbgemm.scala 180:22]
  wire  Gep_24_reset; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_enable_ready; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_enable_valid; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_enable_bits_control; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_Out_0_ready; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_Out_0_valid; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_Out_0_bits_predicate; // @[bbgemm.scala 180:22]
  wire [9:0] Gep_24_io_Out_0_bits_taskID; // @[bbgemm.scala 180:22]
  wire [31:0] Gep_24_io_Out_0_bits_data; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_Out_1_ready; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_Out_1_valid; // @[bbgemm.scala 180:22]
  wire [9:0] Gep_24_io_Out_1_bits_taskID; // @[bbgemm.scala 180:22]
  wire [31:0] Gep_24_io_Out_1_bits_data; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_baseAddress_ready; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_baseAddress_valid; // @[bbgemm.scala 180:22]
  wire [9:0] Gep_24_io_baseAddress_bits_taskID; // @[bbgemm.scala 180:22]
  wire [31:0] Gep_24_io_baseAddress_bits_data; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_idx_0_ready; // @[bbgemm.scala 180:22]
  wire  Gep_24_io_idx_0_valid; // @[bbgemm.scala 180:22]
  wire [31:0] Gep_24_io_idx_0_bits_data; // @[bbgemm.scala 180:22]
  wire  ld_25_clock; // @[bbgemm.scala 183:21]
  wire  ld_25_reset; // @[bbgemm.scala 183:21]
  wire  ld_25_io_enable_ready; // @[bbgemm.scala 183:21]
  wire  ld_25_io_enable_valid; // @[bbgemm.scala 183:21]
  wire [9:0] ld_25_io_enable_bits_taskID; // @[bbgemm.scala 183:21]
  wire  ld_25_io_enable_bits_control; // @[bbgemm.scala 183:21]
  wire  ld_25_io_Out_0_ready; // @[bbgemm.scala 183:21]
  wire  ld_25_io_Out_0_valid; // @[bbgemm.scala 183:21]
  wire [9:0] ld_25_io_Out_0_bits_taskID; // @[bbgemm.scala 183:21]
  wire [31:0] ld_25_io_Out_0_bits_data; // @[bbgemm.scala 183:21]
  wire  ld_25_io_GepAddr_ready; // @[bbgemm.scala 183:21]
  wire  ld_25_io_GepAddr_valid; // @[bbgemm.scala 183:21]
  wire  ld_25_io_GepAddr_bits_predicate; // @[bbgemm.scala 183:21]
  wire [9:0] ld_25_io_GepAddr_bits_taskID; // @[bbgemm.scala 183:21]
  wire [31:0] ld_25_io_GepAddr_bits_data; // @[bbgemm.scala 183:21]
  wire  ld_25_io_memReq_ready; // @[bbgemm.scala 183:21]
  wire  ld_25_io_memReq_valid; // @[bbgemm.scala 183:21]
  wire [31:0] ld_25_io_memReq_bits_address; // @[bbgemm.scala 183:21]
  wire [9:0] ld_25_io_memReq_bits_taskID; // @[bbgemm.scala 183:21]
  wire  ld_25_io_memResp_valid; // @[bbgemm.scala 183:21]
  wire [31:0] ld_25_io_memResp_data; // @[bbgemm.scala 183:21]
  wire  FP_26_clock; // @[bbgemm.scala 187:21]
  wire  FP_26_reset; // @[bbgemm.scala 187:21]
  wire  FP_26_io_enable_ready; // @[bbgemm.scala 187:21]
  wire  FP_26_io_enable_valid; // @[bbgemm.scala 187:21]
  wire [9:0] FP_26_io_enable_bits_taskID; // @[bbgemm.scala 187:21]
  wire  FP_26_io_enable_bits_control; // @[bbgemm.scala 187:21]
  wire  FP_26_io_Out_0_ready; // @[bbgemm.scala 187:21]
  wire  FP_26_io_Out_0_valid; // @[bbgemm.scala 187:21]
  wire [9:0] FP_26_io_Out_0_bits_taskID; // @[bbgemm.scala 187:21]
  wire [31:0] FP_26_io_Out_0_bits_data; // @[bbgemm.scala 187:21]
  wire  FP_26_io_LeftIO_ready; // @[bbgemm.scala 187:21]
  wire  FP_26_io_LeftIO_valid; // @[bbgemm.scala 187:21]
  wire [9:0] FP_26_io_LeftIO_bits_taskID; // @[bbgemm.scala 187:21]
  wire [31:0] FP_26_io_LeftIO_bits_data; // @[bbgemm.scala 187:21]
  wire  FP_26_io_RightIO_ready; // @[bbgemm.scala 187:21]
  wire  FP_26_io_RightIO_valid; // @[bbgemm.scala 187:21]
  wire [9:0] FP_26_io_RightIO_bits_taskID; // @[bbgemm.scala 187:21]
  wire [31:0] FP_26_io_RightIO_bits_data; // @[bbgemm.scala 187:21]
  wire  st_27_clock; // @[bbgemm.scala 190:21]
  wire  st_27_reset; // @[bbgemm.scala 190:21]
  wire  st_27_io_enable_ready; // @[bbgemm.scala 190:21]
  wire  st_27_io_enable_valid; // @[bbgemm.scala 190:21]
  wire [9:0] st_27_io_enable_bits_taskID; // @[bbgemm.scala 190:21]
  wire  st_27_io_enable_bits_control; // @[bbgemm.scala 190:21]
  wire  st_27_io_GepAddr_ready; // @[bbgemm.scala 190:21]
  wire  st_27_io_GepAddr_valid; // @[bbgemm.scala 190:21]
  wire [9:0] st_27_io_GepAddr_bits_taskID; // @[bbgemm.scala 190:21]
  wire [31:0] st_27_io_GepAddr_bits_data; // @[bbgemm.scala 190:21]
  wire  st_27_io_inData_ready; // @[bbgemm.scala 190:21]
  wire  st_27_io_inData_valid; // @[bbgemm.scala 190:21]
  wire [9:0] st_27_io_inData_bits_taskID; // @[bbgemm.scala 190:21]
  wire [31:0] st_27_io_inData_bits_data; // @[bbgemm.scala 190:21]
  wire  st_27_io_memReq_ready; // @[bbgemm.scala 190:21]
  wire  st_27_io_memReq_valid; // @[bbgemm.scala 190:21]
  wire [21:0] st_27_io_memReq_bits_address; // @[bbgemm.scala 190:21]
  wire [31:0] st_27_io_memReq_bits_data; // @[bbgemm.scala 190:21]
  wire [9:0] st_27_io_memReq_bits_taskID; // @[bbgemm.scala 190:21]
  wire  st_27_io_memResp_valid; // @[bbgemm.scala 190:21]
  wire  binaryOp_28_clock; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_reset; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_enable_ready; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_enable_valid; // @[bbgemm.scala 193:27]
  wire [9:0] binaryOp_28_io_enable_bits_taskID; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_enable_bits_control; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_Out_0_ready; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_Out_0_valid; // @[bbgemm.scala 193:27]
  wire [9:0] binaryOp_28_io_Out_0_bits_taskID; // @[bbgemm.scala 193:27]
  wire [31:0] binaryOp_28_io_Out_0_bits_data; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_Out_1_ready; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_Out_1_valid; // @[bbgemm.scala 193:27]
  wire [9:0] binaryOp_28_io_Out_1_bits_taskID; // @[bbgemm.scala 193:27]
  wire [31:0] binaryOp_28_io_Out_1_bits_data; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_LeftIO_ready; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_LeftIO_valid; // @[bbgemm.scala 193:27]
  wire [9:0] binaryOp_28_io_LeftIO_bits_taskID; // @[bbgemm.scala 193:27]
  wire [31:0] binaryOp_28_io_LeftIO_bits_data; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_RightIO_ready; // @[bbgemm.scala 193:27]
  wire  binaryOp_28_io_RightIO_valid; // @[bbgemm.scala 193:27]
  wire [9:0] binaryOp_28_io_RightIO_bits_taskID; // @[bbgemm.scala 193:27]
  wire  icmp_29_clock; // @[bbgemm.scala 196:23]
  wire  icmp_29_reset; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_enable_ready; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_enable_valid; // @[bbgemm.scala 196:23]
  wire [9:0] icmp_29_io_enable_bits_taskID; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_enable_bits_control; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_Out_0_ready; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_Out_0_valid; // @[bbgemm.scala 196:23]
  wire [9:0] icmp_29_io_Out_0_bits_taskID; // @[bbgemm.scala 196:23]
  wire [31:0] icmp_29_io_Out_0_bits_data; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_LeftIO_ready; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_LeftIO_valid; // @[bbgemm.scala 196:23]
  wire [9:0] icmp_29_io_LeftIO_bits_taskID; // @[bbgemm.scala 196:23]
  wire [31:0] icmp_29_io_LeftIO_bits_data; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_RightIO_ready; // @[bbgemm.scala 196:23]
  wire  icmp_29_io_RightIO_valid; // @[bbgemm.scala 196:23]
  wire [9:0] icmp_29_io_RightIO_bits_taskID; // @[bbgemm.scala 196:23]
  wire  br_30_clock; // @[bbgemm.scala 199:21]
  wire  br_30_reset; // @[bbgemm.scala 199:21]
  wire  br_30_io_enable_ready; // @[bbgemm.scala 199:21]
  wire  br_30_io_enable_valid; // @[bbgemm.scala 199:21]
  wire [9:0] br_30_io_enable_bits_taskID; // @[bbgemm.scala 199:21]
  wire  br_30_io_enable_bits_control; // @[bbgemm.scala 199:21]
  wire  br_30_io_CmpIO_ready; // @[bbgemm.scala 199:21]
  wire  br_30_io_CmpIO_valid; // @[bbgemm.scala 199:21]
  wire [9:0] br_30_io_CmpIO_bits_taskID; // @[bbgemm.scala 199:21]
  wire [31:0] br_30_io_CmpIO_bits_data; // @[bbgemm.scala 199:21]
  wire  br_30_io_TrueOutput_0_ready; // @[bbgemm.scala 199:21]
  wire  br_30_io_TrueOutput_0_valid; // @[bbgemm.scala 199:21]
  wire [9:0] br_30_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 199:21]
  wire  br_30_io_TrueOutput_0_bits_control; // @[bbgemm.scala 199:21]
  wire  br_30_io_FalseOutput_0_ready; // @[bbgemm.scala 199:21]
  wire  br_30_io_FalseOutput_0_valid; // @[bbgemm.scala 199:21]
  wire [9:0] br_30_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 199:21]
  wire  br_30_io_FalseOutput_0_bits_control; // @[bbgemm.scala 199:21]
  wire  binaryOp_31_clock; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_reset; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_enable_ready; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_enable_valid; // @[bbgemm.scala 202:27]
  wire [9:0] binaryOp_31_io_enable_bits_taskID; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_enable_bits_control; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_Out_0_ready; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_Out_0_valid; // @[bbgemm.scala 202:27]
  wire [9:0] binaryOp_31_io_Out_0_bits_taskID; // @[bbgemm.scala 202:27]
  wire [31:0] binaryOp_31_io_Out_0_bits_data; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_Out_1_ready; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_Out_1_valid; // @[bbgemm.scala 202:27]
  wire [9:0] binaryOp_31_io_Out_1_bits_taskID; // @[bbgemm.scala 202:27]
  wire [31:0] binaryOp_31_io_Out_1_bits_data; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_LeftIO_ready; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_LeftIO_valid; // @[bbgemm.scala 202:27]
  wire [9:0] binaryOp_31_io_LeftIO_bits_taskID; // @[bbgemm.scala 202:27]
  wire [31:0] binaryOp_31_io_LeftIO_bits_data; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_RightIO_ready; // @[bbgemm.scala 202:27]
  wire  binaryOp_31_io_RightIO_valid; // @[bbgemm.scala 202:27]
  wire [9:0] binaryOp_31_io_RightIO_bits_taskID; // @[bbgemm.scala 202:27]
  wire  icmp_32_clock; // @[bbgemm.scala 205:23]
  wire  icmp_32_reset; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_enable_ready; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_enable_valid; // @[bbgemm.scala 205:23]
  wire [9:0] icmp_32_io_enable_bits_taskID; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_enable_bits_control; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_Out_0_ready; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_Out_0_valid; // @[bbgemm.scala 205:23]
  wire [9:0] icmp_32_io_Out_0_bits_taskID; // @[bbgemm.scala 205:23]
  wire [31:0] icmp_32_io_Out_0_bits_data; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_LeftIO_ready; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_LeftIO_valid; // @[bbgemm.scala 205:23]
  wire [9:0] icmp_32_io_LeftIO_bits_taskID; // @[bbgemm.scala 205:23]
  wire [31:0] icmp_32_io_LeftIO_bits_data; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_RightIO_ready; // @[bbgemm.scala 205:23]
  wire  icmp_32_io_RightIO_valid; // @[bbgemm.scala 205:23]
  wire [9:0] icmp_32_io_RightIO_bits_taskID; // @[bbgemm.scala 205:23]
  wire  br_33_clock; // @[bbgemm.scala 208:21]
  wire  br_33_reset; // @[bbgemm.scala 208:21]
  wire  br_33_io_enable_ready; // @[bbgemm.scala 208:21]
  wire  br_33_io_enable_valid; // @[bbgemm.scala 208:21]
  wire [9:0] br_33_io_enable_bits_taskID; // @[bbgemm.scala 208:21]
  wire  br_33_io_enable_bits_control; // @[bbgemm.scala 208:21]
  wire  br_33_io_CmpIO_ready; // @[bbgemm.scala 208:21]
  wire  br_33_io_CmpIO_valid; // @[bbgemm.scala 208:21]
  wire [9:0] br_33_io_CmpIO_bits_taskID; // @[bbgemm.scala 208:21]
  wire [31:0] br_33_io_CmpIO_bits_data; // @[bbgemm.scala 208:21]
  wire  br_33_io_TrueOutput_0_ready; // @[bbgemm.scala 208:21]
  wire  br_33_io_TrueOutput_0_valid; // @[bbgemm.scala 208:21]
  wire [9:0] br_33_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 208:21]
  wire  br_33_io_TrueOutput_0_bits_control; // @[bbgemm.scala 208:21]
  wire  br_33_io_FalseOutput_0_ready; // @[bbgemm.scala 208:21]
  wire  br_33_io_FalseOutput_0_valid; // @[bbgemm.scala 208:21]
  wire [9:0] br_33_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 208:21]
  wire  br_33_io_FalseOutput_0_bits_control; // @[bbgemm.scala 208:21]
  wire  binaryOp_34_clock; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_reset; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_enable_ready; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_enable_valid; // @[bbgemm.scala 211:27]
  wire [9:0] binaryOp_34_io_enable_bits_taskID; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_enable_bits_control; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_Out_0_ready; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_Out_0_valid; // @[bbgemm.scala 211:27]
  wire [9:0] binaryOp_34_io_Out_0_bits_taskID; // @[bbgemm.scala 211:27]
  wire [31:0] binaryOp_34_io_Out_0_bits_data; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_Out_1_ready; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_Out_1_valid; // @[bbgemm.scala 211:27]
  wire [9:0] binaryOp_34_io_Out_1_bits_taskID; // @[bbgemm.scala 211:27]
  wire [31:0] binaryOp_34_io_Out_1_bits_data; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_LeftIO_ready; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_LeftIO_valid; // @[bbgemm.scala 211:27]
  wire [9:0] binaryOp_34_io_LeftIO_bits_taskID; // @[bbgemm.scala 211:27]
  wire [31:0] binaryOp_34_io_LeftIO_bits_data; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_RightIO_ready; // @[bbgemm.scala 211:27]
  wire  binaryOp_34_io_RightIO_valid; // @[bbgemm.scala 211:27]
  wire [9:0] binaryOp_34_io_RightIO_bits_taskID; // @[bbgemm.scala 211:27]
  wire  icmp_35_clock; // @[bbgemm.scala 214:23]
  wire  icmp_35_reset; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_enable_ready; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_enable_valid; // @[bbgemm.scala 214:23]
  wire [9:0] icmp_35_io_enable_bits_taskID; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_enable_bits_control; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_Out_0_ready; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_Out_0_valid; // @[bbgemm.scala 214:23]
  wire [9:0] icmp_35_io_Out_0_bits_taskID; // @[bbgemm.scala 214:23]
  wire [31:0] icmp_35_io_Out_0_bits_data; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_LeftIO_ready; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_LeftIO_valid; // @[bbgemm.scala 214:23]
  wire [9:0] icmp_35_io_LeftIO_bits_taskID; // @[bbgemm.scala 214:23]
  wire [31:0] icmp_35_io_LeftIO_bits_data; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_RightIO_ready; // @[bbgemm.scala 214:23]
  wire  icmp_35_io_RightIO_valid; // @[bbgemm.scala 214:23]
  wire [9:0] icmp_35_io_RightIO_bits_taskID; // @[bbgemm.scala 214:23]
  wire  br_36_clock; // @[bbgemm.scala 217:21]
  wire  br_36_reset; // @[bbgemm.scala 217:21]
  wire  br_36_io_enable_ready; // @[bbgemm.scala 217:21]
  wire  br_36_io_enable_valid; // @[bbgemm.scala 217:21]
  wire [9:0] br_36_io_enable_bits_taskID; // @[bbgemm.scala 217:21]
  wire  br_36_io_enable_bits_control; // @[bbgemm.scala 217:21]
  wire  br_36_io_CmpIO_ready; // @[bbgemm.scala 217:21]
  wire  br_36_io_CmpIO_valid; // @[bbgemm.scala 217:21]
  wire [9:0] br_36_io_CmpIO_bits_taskID; // @[bbgemm.scala 217:21]
  wire [31:0] br_36_io_CmpIO_bits_data; // @[bbgemm.scala 217:21]
  wire  br_36_io_TrueOutput_0_ready; // @[bbgemm.scala 217:21]
  wire  br_36_io_TrueOutput_0_valid; // @[bbgemm.scala 217:21]
  wire [9:0] br_36_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 217:21]
  wire  br_36_io_TrueOutput_0_bits_control; // @[bbgemm.scala 217:21]
  wire  br_36_io_FalseOutput_0_ready; // @[bbgemm.scala 217:21]
  wire  br_36_io_FalseOutput_0_valid; // @[bbgemm.scala 217:21]
  wire [9:0] br_36_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 217:21]
  wire  br_36_io_FalseOutput_0_bits_control; // @[bbgemm.scala 217:21]
  wire  binaryOp_37_clock; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_reset; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_enable_ready; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_enable_valid; // @[bbgemm.scala 220:27]
  wire [9:0] binaryOp_37_io_enable_bits_taskID; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_enable_bits_control; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_Out_0_ready; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_Out_0_valid; // @[bbgemm.scala 220:27]
  wire [9:0] binaryOp_37_io_Out_0_bits_taskID; // @[bbgemm.scala 220:27]
  wire [31:0] binaryOp_37_io_Out_0_bits_data; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_Out_1_ready; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_Out_1_valid; // @[bbgemm.scala 220:27]
  wire [9:0] binaryOp_37_io_Out_1_bits_taskID; // @[bbgemm.scala 220:27]
  wire [31:0] binaryOp_37_io_Out_1_bits_data; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_LeftIO_ready; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_LeftIO_valid; // @[bbgemm.scala 220:27]
  wire [9:0] binaryOp_37_io_LeftIO_bits_taskID; // @[bbgemm.scala 220:27]
  wire [31:0] binaryOp_37_io_LeftIO_bits_data; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_RightIO_ready; // @[bbgemm.scala 220:27]
  wire  binaryOp_37_io_RightIO_valid; // @[bbgemm.scala 220:27]
  wire [9:0] binaryOp_37_io_RightIO_bits_taskID; // @[bbgemm.scala 220:27]
  wire  icmp_38_clock; // @[bbgemm.scala 223:23]
  wire  icmp_38_reset; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_enable_ready; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_enable_valid; // @[bbgemm.scala 223:23]
  wire [9:0] icmp_38_io_enable_bits_taskID; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_enable_bits_control; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_Out_0_ready; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_Out_0_valid; // @[bbgemm.scala 223:23]
  wire [9:0] icmp_38_io_Out_0_bits_taskID; // @[bbgemm.scala 223:23]
  wire [31:0] icmp_38_io_Out_0_bits_data; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_LeftIO_ready; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_LeftIO_valid; // @[bbgemm.scala 223:23]
  wire [9:0] icmp_38_io_LeftIO_bits_taskID; // @[bbgemm.scala 223:23]
  wire [31:0] icmp_38_io_LeftIO_bits_data; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_RightIO_ready; // @[bbgemm.scala 223:23]
  wire  icmp_38_io_RightIO_valid; // @[bbgemm.scala 223:23]
  wire [9:0] icmp_38_io_RightIO_bits_taskID; // @[bbgemm.scala 223:23]
  wire  br_39_clock; // @[bbgemm.scala 226:21]
  wire  br_39_reset; // @[bbgemm.scala 226:21]
  wire  br_39_io_enable_ready; // @[bbgemm.scala 226:21]
  wire  br_39_io_enable_valid; // @[bbgemm.scala 226:21]
  wire [9:0] br_39_io_enable_bits_taskID; // @[bbgemm.scala 226:21]
  wire  br_39_io_enable_bits_control; // @[bbgemm.scala 226:21]
  wire  br_39_io_CmpIO_ready; // @[bbgemm.scala 226:21]
  wire  br_39_io_CmpIO_valid; // @[bbgemm.scala 226:21]
  wire [9:0] br_39_io_CmpIO_bits_taskID; // @[bbgemm.scala 226:21]
  wire [31:0] br_39_io_CmpIO_bits_data; // @[bbgemm.scala 226:21]
  wire  br_39_io_TrueOutput_0_ready; // @[bbgemm.scala 226:21]
  wire  br_39_io_TrueOutput_0_valid; // @[bbgemm.scala 226:21]
  wire [9:0] br_39_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 226:21]
  wire  br_39_io_TrueOutput_0_bits_control; // @[bbgemm.scala 226:21]
  wire  br_39_io_FalseOutput_0_ready; // @[bbgemm.scala 226:21]
  wire  br_39_io_FalseOutput_0_valid; // @[bbgemm.scala 226:21]
  wire [9:0] br_39_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 226:21]
  wire  br_39_io_FalseOutput_0_bits_control; // @[bbgemm.scala 226:21]
  wire  binaryOp_40_clock; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_reset; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_enable_ready; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_enable_valid; // @[bbgemm.scala 229:27]
  wire [9:0] binaryOp_40_io_enable_bits_taskID; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_enable_bits_control; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_Out_0_ready; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_Out_0_valid; // @[bbgemm.scala 229:27]
  wire [9:0] binaryOp_40_io_Out_0_bits_taskID; // @[bbgemm.scala 229:27]
  wire [31:0] binaryOp_40_io_Out_0_bits_data; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_Out_1_ready; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_Out_1_valid; // @[bbgemm.scala 229:27]
  wire [9:0] binaryOp_40_io_Out_1_bits_taskID; // @[bbgemm.scala 229:27]
  wire [31:0] binaryOp_40_io_Out_1_bits_data; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_LeftIO_ready; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_LeftIO_valid; // @[bbgemm.scala 229:27]
  wire [9:0] binaryOp_40_io_LeftIO_bits_taskID; // @[bbgemm.scala 229:27]
  wire [31:0] binaryOp_40_io_LeftIO_bits_data; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_RightIO_ready; // @[bbgemm.scala 229:27]
  wire  binaryOp_40_io_RightIO_valid; // @[bbgemm.scala 229:27]
  wire [9:0] binaryOp_40_io_RightIO_bits_taskID; // @[bbgemm.scala 229:27]
  wire  icmp_41_clock; // @[bbgemm.scala 232:23]
  wire  icmp_41_reset; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_enable_ready; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_enable_valid; // @[bbgemm.scala 232:23]
  wire [9:0] icmp_41_io_enable_bits_taskID; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_enable_bits_control; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_Out_0_ready; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_Out_0_valid; // @[bbgemm.scala 232:23]
  wire [9:0] icmp_41_io_Out_0_bits_taskID; // @[bbgemm.scala 232:23]
  wire [31:0] icmp_41_io_Out_0_bits_data; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_LeftIO_ready; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_LeftIO_valid; // @[bbgemm.scala 232:23]
  wire [9:0] icmp_41_io_LeftIO_bits_taskID; // @[bbgemm.scala 232:23]
  wire [31:0] icmp_41_io_LeftIO_bits_data; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_RightIO_ready; // @[bbgemm.scala 232:23]
  wire  icmp_41_io_RightIO_valid; // @[bbgemm.scala 232:23]
  wire [9:0] icmp_41_io_RightIO_bits_taskID; // @[bbgemm.scala 232:23]
  wire  br_42_clock; // @[bbgemm.scala 235:21]
  wire  br_42_reset; // @[bbgemm.scala 235:21]
  wire  br_42_io_enable_ready; // @[bbgemm.scala 235:21]
  wire  br_42_io_enable_valid; // @[bbgemm.scala 235:21]
  wire [9:0] br_42_io_enable_bits_taskID; // @[bbgemm.scala 235:21]
  wire  br_42_io_enable_bits_control; // @[bbgemm.scala 235:21]
  wire  br_42_io_CmpIO_ready; // @[bbgemm.scala 235:21]
  wire  br_42_io_CmpIO_valid; // @[bbgemm.scala 235:21]
  wire [9:0] br_42_io_CmpIO_bits_taskID; // @[bbgemm.scala 235:21]
  wire [31:0] br_42_io_CmpIO_bits_data; // @[bbgemm.scala 235:21]
  wire  br_42_io_TrueOutput_0_ready; // @[bbgemm.scala 235:21]
  wire  br_42_io_TrueOutput_0_valid; // @[bbgemm.scala 235:21]
  wire [9:0] br_42_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 235:21]
  wire  br_42_io_TrueOutput_0_bits_control; // @[bbgemm.scala 235:21]
  wire  br_42_io_FalseOutput_0_ready; // @[bbgemm.scala 235:21]
  wire  br_42_io_FalseOutput_0_valid; // @[bbgemm.scala 235:21]
  wire [9:0] br_42_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 235:21]
  wire  br_42_io_FalseOutput_0_bits_control; // @[bbgemm.scala 235:21]
  wire  ret_43_clock; // @[bbgemm.scala 238:22]
  wire  ret_43_reset; // @[bbgemm.scala 238:22]
  wire  ret_43_io_In_enable_ready; // @[bbgemm.scala 238:22]
  wire  ret_43_io_In_enable_valid; // @[bbgemm.scala 238:22]
  wire [9:0] ret_43_io_In_enable_bits_taskID; // @[bbgemm.scala 238:22]
  wire  ret_43_io_In_enable_bits_control; // @[bbgemm.scala 238:22]
  wire  ret_43_io_Out_ready; // @[bbgemm.scala 238:22]
  wire  ret_43_io_Out_valid; // @[bbgemm.scala 238:22]
  wire [9:0] ret_43_io_Out_bits_enable_taskID; // @[bbgemm.scala 238:22]
  wire  ret_43_io_Out_bits_enable_control; // @[bbgemm.scala 238:22]
  wire  const0_clock; // @[bbgemm.scala 247:22]
  wire  const0_reset; // @[bbgemm.scala 247:22]
  wire  const0_io_enable_ready; // @[bbgemm.scala 247:22]
  wire  const0_io_enable_valid; // @[bbgemm.scala 247:22]
  wire [9:0] const0_io_enable_bits_taskID; // @[bbgemm.scala 247:22]
  wire  const0_io_Out_ready; // @[bbgemm.scala 247:22]
  wire  const0_io_Out_valid; // @[bbgemm.scala 247:22]
  wire [9:0] const0_io_Out_bits_taskID; // @[bbgemm.scala 247:22]
  wire  const1_clock; // @[bbgemm.scala 250:22]
  wire  const1_reset; // @[bbgemm.scala 250:22]
  wire  const1_io_enable_ready; // @[bbgemm.scala 250:22]
  wire  const1_io_enable_valid; // @[bbgemm.scala 250:22]
  wire [9:0] const1_io_enable_bits_taskID; // @[bbgemm.scala 250:22]
  wire  const1_io_Out_ready; // @[bbgemm.scala 250:22]
  wire  const1_io_Out_valid; // @[bbgemm.scala 250:22]
  wire [9:0] const1_io_Out_bits_taskID; // @[bbgemm.scala 250:22]
  wire  const2_clock; // @[bbgemm.scala 253:22]
  wire  const2_reset; // @[bbgemm.scala 253:22]
  wire  const2_io_enable_ready; // @[bbgemm.scala 253:22]
  wire  const2_io_enable_valid; // @[bbgemm.scala 253:22]
  wire [9:0] const2_io_enable_bits_taskID; // @[bbgemm.scala 253:22]
  wire  const2_io_Out_ready; // @[bbgemm.scala 253:22]
  wire  const2_io_Out_valid; // @[bbgemm.scala 253:22]
  wire [9:0] const2_io_Out_bits_taskID; // @[bbgemm.scala 253:22]
  wire  const3_clock; // @[bbgemm.scala 256:22]
  wire  const3_reset; // @[bbgemm.scala 256:22]
  wire  const3_io_enable_ready; // @[bbgemm.scala 256:22]
  wire  const3_io_enable_valid; // @[bbgemm.scala 256:22]
  wire  const3_io_Out_ready; // @[bbgemm.scala 256:22]
  wire  const3_io_Out_valid; // @[bbgemm.scala 256:22]
  wire  const4_clock; // @[bbgemm.scala 259:22]
  wire  const4_reset; // @[bbgemm.scala 259:22]
  wire  const4_io_enable_ready; // @[bbgemm.scala 259:22]
  wire  const4_io_enable_valid; // @[bbgemm.scala 259:22]
  wire [9:0] const4_io_enable_bits_taskID; // @[bbgemm.scala 259:22]
  wire  const4_io_Out_ready; // @[bbgemm.scala 259:22]
  wire  const4_io_Out_valid; // @[bbgemm.scala 259:22]
  wire [9:0] const4_io_Out_bits_taskID; // @[bbgemm.scala 259:22]
  wire  const5_clock; // @[bbgemm.scala 262:22]
  wire  const5_reset; // @[bbgemm.scala 262:22]
  wire  const5_io_enable_ready; // @[bbgemm.scala 262:22]
  wire  const5_io_enable_valid; // @[bbgemm.scala 262:22]
  wire  const5_io_Out_ready; // @[bbgemm.scala 262:22]
  wire  const5_io_Out_valid; // @[bbgemm.scala 262:22]
  wire  const6_clock; // @[bbgemm.scala 265:22]
  wire  const6_reset; // @[bbgemm.scala 265:22]
  wire  const6_io_enable_ready; // @[bbgemm.scala 265:22]
  wire  const6_io_enable_valid; // @[bbgemm.scala 265:22]
  wire [9:0] const6_io_enable_bits_taskID; // @[bbgemm.scala 265:22]
  wire  const6_io_Out_ready; // @[bbgemm.scala 265:22]
  wire  const6_io_Out_valid; // @[bbgemm.scala 265:22]
  wire [9:0] const6_io_Out_bits_taskID; // @[bbgemm.scala 265:22]
  wire  const7_clock; // @[bbgemm.scala 268:22]
  wire  const7_reset; // @[bbgemm.scala 268:22]
  wire  const7_io_enable_ready; // @[bbgemm.scala 268:22]
  wire  const7_io_enable_valid; // @[bbgemm.scala 268:22]
  wire [9:0] const7_io_enable_bits_taskID; // @[bbgemm.scala 268:22]
  wire  const7_io_Out_ready; // @[bbgemm.scala 268:22]
  wire  const7_io_Out_valid; // @[bbgemm.scala 268:22]
  wire [9:0] const7_io_Out_bits_taskID; // @[bbgemm.scala 268:22]
  wire  const8_clock; // @[bbgemm.scala 271:22]
  wire  const8_reset; // @[bbgemm.scala 271:22]
  wire  const8_io_enable_ready; // @[bbgemm.scala 271:22]
  wire  const8_io_enable_valid; // @[bbgemm.scala 271:22]
  wire [9:0] const8_io_enable_bits_taskID; // @[bbgemm.scala 271:22]
  wire  const8_io_Out_ready; // @[bbgemm.scala 271:22]
  wire  const8_io_Out_valid; // @[bbgemm.scala 271:22]
  wire [9:0] const8_io_Out_bits_taskID; // @[bbgemm.scala 271:22]
  wire  const9_clock; // @[bbgemm.scala 274:22]
  wire  const9_reset; // @[bbgemm.scala 274:22]
  wire  const9_io_enable_ready; // @[bbgemm.scala 274:22]
  wire  const9_io_enable_valid; // @[bbgemm.scala 274:22]
  wire [9:0] const9_io_enable_bits_taskID; // @[bbgemm.scala 274:22]
  wire  const9_io_Out_ready; // @[bbgemm.scala 274:22]
  wire  const9_io_Out_valid; // @[bbgemm.scala 274:22]
  wire [9:0] const9_io_Out_bits_taskID; // @[bbgemm.scala 274:22]
  wire  const10_clock; // @[bbgemm.scala 277:23]
  wire  const10_reset; // @[bbgemm.scala 277:23]
  wire  const10_io_enable_ready; // @[bbgemm.scala 277:23]
  wire  const10_io_enable_valid; // @[bbgemm.scala 277:23]
  wire [9:0] const10_io_enable_bits_taskID; // @[bbgemm.scala 277:23]
  wire  const10_io_Out_ready; // @[bbgemm.scala 277:23]
  wire  const10_io_Out_valid; // @[bbgemm.scala 277:23]
  wire [9:0] const10_io_Out_bits_taskID; // @[bbgemm.scala 277:23]
  wire  const11_clock; // @[bbgemm.scala 280:23]
  wire  const11_reset; // @[bbgemm.scala 280:23]
  wire  const11_io_enable_ready; // @[bbgemm.scala 280:23]
  wire  const11_io_enable_valid; // @[bbgemm.scala 280:23]
  wire [9:0] const11_io_enable_bits_taskID; // @[bbgemm.scala 280:23]
  wire  const11_io_Out_ready; // @[bbgemm.scala 280:23]
  wire  const11_io_Out_valid; // @[bbgemm.scala 280:23]
  wire [9:0] const11_io_Out_bits_taskID; // @[bbgemm.scala 280:23]
  wire  const12_clock; // @[bbgemm.scala 283:23]
  wire  const12_reset; // @[bbgemm.scala 283:23]
  wire  const12_io_enable_ready; // @[bbgemm.scala 283:23]
  wire  const12_io_enable_valid; // @[bbgemm.scala 283:23]
  wire [9:0] const12_io_enable_bits_taskID; // @[bbgemm.scala 283:23]
  wire  const12_io_Out_ready; // @[bbgemm.scala 283:23]
  wire  const12_io_Out_valid; // @[bbgemm.scala 283:23]
  wire [9:0] const12_io_Out_bits_taskID; // @[bbgemm.scala 283:23]
  wire  const13_clock; // @[bbgemm.scala 286:23]
  wire  const13_reset; // @[bbgemm.scala 286:23]
  wire  const13_io_enable_ready; // @[bbgemm.scala 286:23]
  wire  const13_io_enable_valid; // @[bbgemm.scala 286:23]
  wire [9:0] const13_io_enable_bits_taskID; // @[bbgemm.scala 286:23]
  wire  const13_io_Out_ready; // @[bbgemm.scala 286:23]
  wire  const13_io_Out_valid; // @[bbgemm.scala 286:23]
  wire [9:0] const13_io_Out_bits_taskID; // @[bbgemm.scala 286:23]
  wire  const14_clock; // @[bbgemm.scala 289:23]
  wire  const14_reset; // @[bbgemm.scala 289:23]
  wire  const14_io_enable_ready; // @[bbgemm.scala 289:23]
  wire  const14_io_enable_valid; // @[bbgemm.scala 289:23]
  wire [9:0] const14_io_enable_bits_taskID; // @[bbgemm.scala 289:23]
  wire  const14_io_Out_ready; // @[bbgemm.scala 289:23]
  wire  const14_io_Out_valid; // @[bbgemm.scala 289:23]
  wire [9:0] const14_io_Out_bits_taskID; // @[bbgemm.scala 289:23]
  wire  const15_clock; // @[bbgemm.scala 292:23]
  wire  const15_reset; // @[bbgemm.scala 292:23]
  wire  const15_io_enable_ready; // @[bbgemm.scala 292:23]
  wire  const15_io_enable_valid; // @[bbgemm.scala 292:23]
  wire [9:0] const15_io_enable_bits_taskID; // @[bbgemm.scala 292:23]
  wire  const15_io_Out_ready; // @[bbgemm.scala 292:23]
  wire  const15_io_Out_valid; // @[bbgemm.scala 292:23]
  wire [9:0] const15_io_Out_bits_taskID; // @[bbgemm.scala 292:23]
  wire  const16_clock; // @[bbgemm.scala 295:23]
  wire  const16_reset; // @[bbgemm.scala 295:23]
  wire  const16_io_enable_ready; // @[bbgemm.scala 295:23]
  wire  const16_io_enable_valid; // @[bbgemm.scala 295:23]
  wire [9:0] const16_io_enable_bits_taskID; // @[bbgemm.scala 295:23]
  wire  const16_io_Out_ready; // @[bbgemm.scala 295:23]
  wire  const16_io_Out_valid; // @[bbgemm.scala 295:23]
  wire [9:0] const16_io_Out_bits_taskID; // @[bbgemm.scala 295:23]
  UnifiedController MemCtrl ( // @[bbgemm.scala 45:23]
    .clock(MemCtrl_clock),
    .reset(MemCtrl_reset),
    .io_WriteIn_0_ready(MemCtrl_io_WriteIn_0_ready),
    .io_WriteIn_0_valid(MemCtrl_io_WriteIn_0_valid),
    .io_WriteIn_0_bits_address(MemCtrl_io_WriteIn_0_bits_address),
    .io_WriteIn_0_bits_data(MemCtrl_io_WriteIn_0_bits_data),
    .io_WriteIn_0_bits_taskID(MemCtrl_io_WriteIn_0_bits_taskID),
    .io_WriteOut_0_valid(MemCtrl_io_WriteOut_0_valid),
    .io_ReadIn_0_ready(MemCtrl_io_ReadIn_0_ready),
    .io_ReadIn_0_valid(MemCtrl_io_ReadIn_0_valid),
    .io_ReadIn_0_bits_address(MemCtrl_io_ReadIn_0_bits_address),
    .io_ReadIn_0_bits_taskID(MemCtrl_io_ReadIn_0_bits_taskID),
    .io_ReadIn_1_ready(MemCtrl_io_ReadIn_1_ready),
    .io_ReadIn_1_valid(MemCtrl_io_ReadIn_1_valid),
    .io_ReadIn_1_bits_address(MemCtrl_io_ReadIn_1_bits_address),
    .io_ReadIn_1_bits_taskID(MemCtrl_io_ReadIn_1_bits_taskID),
    .io_ReadIn_2_ready(MemCtrl_io_ReadIn_2_ready),
    .io_ReadIn_2_valid(MemCtrl_io_ReadIn_2_valid),
    .io_ReadIn_2_bits_address(MemCtrl_io_ReadIn_2_bits_address),
    .io_ReadIn_2_bits_taskID(MemCtrl_io_ReadIn_2_bits_taskID),
    .io_ReadOut_0_valid(MemCtrl_io_ReadOut_0_valid),
    .io_ReadOut_0_data(MemCtrl_io_ReadOut_0_data),
    .io_ReadOut_1_valid(MemCtrl_io_ReadOut_1_valid),
    .io_ReadOut_1_data(MemCtrl_io_ReadOut_1_data),
    .io_ReadOut_2_valid(MemCtrl_io_ReadOut_2_valid),
    .io_ReadOut_2_data(MemCtrl_io_ReadOut_2_data),
    .io_MemResp_valid(MemCtrl_io_MemResp_valid),
    .io_MemResp_bits_data(MemCtrl_io_MemResp_bits_data),
    .io_MemResp_bits_tag(MemCtrl_io_MemResp_bits_tag),
    .io_MemResp_bits_iswrite(MemCtrl_io_MemResp_bits_iswrite),
    .io_MemReq_ready(MemCtrl_io_MemReq_ready),
    .io_MemReq_valid(MemCtrl_io_MemReq_valid),
    .io_MemReq_bits_addr(MemCtrl_io_MemReq_bits_addr),
    .io_MemReq_bits_data(MemCtrl_io_MemReq_bits_data),
    .io_MemReq_bits_mask(MemCtrl_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(MemCtrl_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(MemCtrl_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(MemCtrl_io_MemReq_bits_iswrite)
  );
  SplitCallNew InputSplitter ( // @[bbgemm.scala 53:29]
    .clock(InputSplitter_clock),
    .reset(InputSplitter_reset),
    .io_In_ready(InputSplitter_io_In_ready),
    .io_In_valid(InputSplitter_io_In_valid),
    .io_In_bits_enable_taskID(InputSplitter_io_In_bits_enable_taskID),
    .io_In_bits_enable_control(InputSplitter_io_In_bits_enable_control),
    .io_In_bits_data_field2_taskID(InputSplitter_io_In_bits_data_field2_taskID),
    .io_In_bits_data_field2_data(InputSplitter_io_In_bits_data_field2_data),
    .io_In_bits_data_field1_taskID(InputSplitter_io_In_bits_data_field1_taskID),
    .io_In_bits_data_field1_data(InputSplitter_io_In_bits_data_field1_data),
    .io_In_bits_data_field0_taskID(InputSplitter_io_In_bits_data_field0_taskID),
    .io_In_bits_data_field0_data(InputSplitter_io_In_bits_data_field0_data),
    .io_Out_enable_ready(InputSplitter_io_Out_enable_ready),
    .io_Out_enable_valid(InputSplitter_io_Out_enable_valid),
    .io_Out_enable_bits_taskID(InputSplitter_io_Out_enable_bits_taskID),
    .io_Out_enable_bits_control(InputSplitter_io_Out_enable_bits_control),
    .io_Out_data_field2_0_ready(InputSplitter_io_Out_data_field2_0_ready),
    .io_Out_data_field2_0_valid(InputSplitter_io_Out_data_field2_0_valid),
    .io_Out_data_field2_0_bits_taskID(InputSplitter_io_Out_data_field2_0_bits_taskID),
    .io_Out_data_field2_0_bits_data(InputSplitter_io_Out_data_field2_0_bits_data),
    .io_Out_data_field1_0_ready(InputSplitter_io_Out_data_field1_0_ready),
    .io_Out_data_field1_0_valid(InputSplitter_io_Out_data_field1_0_valid),
    .io_Out_data_field1_0_bits_taskID(InputSplitter_io_Out_data_field1_0_bits_taskID),
    .io_Out_data_field1_0_bits_data(InputSplitter_io_Out_data_field1_0_bits_data),
    .io_Out_data_field0_0_ready(InputSplitter_io_Out_data_field0_0_ready),
    .io_Out_data_field0_0_valid(InputSplitter_io_Out_data_field0_0_valid),
    .io_Out_data_field0_0_bits_taskID(InputSplitter_io_Out_data_field0_0_bits_taskID),
    .io_Out_data_field0_0_bits_data(InputSplitter_io_Out_data_field0_0_bits_data)
  );
  LoopBlockNode Loop_0 ( // @[bbgemm.scala 62:22]
    .clock(Loop_0_clock),
    .reset(Loop_0_reset),
    .io_enable_ready(Loop_0_io_enable_ready),
    .io_enable_valid(Loop_0_io_enable_valid),
    .io_enable_bits_taskID(Loop_0_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_0_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_0_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_0_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_0_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_0_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_0_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_taskID(Loop_0_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_0_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_0_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_0_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_0_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_0_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_0_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_taskID(Loop_0_io_InLiveIn_3_bits_taskID),
    .io_InLiveIn_3_bits_data(Loop_0_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_0_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_0_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_taskID(Loop_0_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_0_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_0_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_0_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_0_io_InLiveIn_5_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_0_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_0_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_0_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field5_1_ready(Loop_0_io_OutLiveIn_field5_1_ready),
    .io_OutLiveIn_field5_1_valid(Loop_0_io_OutLiveIn_field5_1_valid),
    .io_OutLiveIn_field5_1_bits_data(Loop_0_io_OutLiveIn_field5_1_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_0_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_0_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_0_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_0_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_0_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_0_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_taskID(Loop_0_io_OutLiveIn_field3_0_bits_taskID),
    .io_OutLiveIn_field3_0_bits_data(Loop_0_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_0_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_0_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_0_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_0_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_0_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_0_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_0_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_0_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_0_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_0_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_0_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_0_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_0_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_0_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_0_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_0_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_0_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_0_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_0_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_0_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_0_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_0_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_0_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_0_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_0_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_0_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_0_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_0_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_0_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_0_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_0_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_0_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_0_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_0_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_0_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_0_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_0_io_loopExit_0_bits_control)
  );
  LoopBlockNode_1 Loop_1 ( // @[bbgemm.scala 64:22]
    .clock(Loop_1_clock),
    .reset(Loop_1_reset),
    .io_enable_ready(Loop_1_io_enable_ready),
    .io_enable_valid(Loop_1_io_enable_valid),
    .io_enable_bits_taskID(Loop_1_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_1_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_1_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_1_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_1_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_1_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_1_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_taskID(Loop_1_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_1_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_1_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_1_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_1_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_1_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_1_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_1_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_1_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_1_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_1_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_data(Loop_1_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_1_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_1_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_taskID(Loop_1_io_InLiveIn_5_bits_taskID),
    .io_InLiveIn_5_bits_data(Loop_1_io_InLiveIn_5_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_1_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_1_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_taskID(Loop_1_io_OutLiveIn_field5_0_bits_taskID),
    .io_OutLiveIn_field5_0_bits_data(Loop_1_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_1_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_1_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_data(Loop_1_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field4_1_ready(Loop_1_io_OutLiveIn_field4_1_ready),
    .io_OutLiveIn_field4_1_valid(Loop_1_io_OutLiveIn_field4_1_valid),
    .io_OutLiveIn_field4_1_bits_data(Loop_1_io_OutLiveIn_field4_1_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_1_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_1_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_1_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_1_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_1_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_1_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_1_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_1_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_1_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_1_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_1_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_1_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_1_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_1_io_OutLiveIn_field0_0_bits_data),
    .io_OutLiveIn_field0_1_ready(Loop_1_io_OutLiveIn_field0_1_ready),
    .io_OutLiveIn_field0_1_valid(Loop_1_io_OutLiveIn_field0_1_valid),
    .io_OutLiveIn_field0_1_bits_data(Loop_1_io_OutLiveIn_field0_1_bits_data),
    .io_activate_loop_start_ready(Loop_1_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_1_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_1_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_1_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_1_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_1_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_1_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_1_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_1_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_1_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_1_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_1_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_1_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_1_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_1_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_1_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_1_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_1_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_1_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_1_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_1_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_1_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_1_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_1_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_1_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_1_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_1_io_loopExit_0_bits_control)
  );
  LoopBlockNode_2 Loop_2 ( // @[bbgemm.scala 66:22]
    .clock(Loop_2_clock),
    .reset(Loop_2_reset),
    .io_enable_ready(Loop_2_io_enable_ready),
    .io_enable_valid(Loop_2_io_enable_valid),
    .io_enable_bits_taskID(Loop_2_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_2_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_2_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_2_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_2_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_2_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_2_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_taskID(Loop_2_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_2_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_2_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_2_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_2_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_2_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_2_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_2_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_taskID(Loop_2_io_InLiveIn_3_bits_taskID),
    .io_InLiveIn_3_bits_data(Loop_2_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_2_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_2_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_data(Loop_2_io_InLiveIn_4_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_2_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_2_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_data(Loop_2_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_2_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_2_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_taskID(Loop_2_io_OutLiveIn_field3_0_bits_taskID),
    .io_OutLiveIn_field3_0_bits_data(Loop_2_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_2_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_2_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_2_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_2_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_2_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_2_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_2_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_2_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_2_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_2_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_2_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_2_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_2_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_2_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_2_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_2_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_2_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_2_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_2_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_2_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_2_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_2_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_2_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_2_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_2_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_2_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_2_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_2_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_2_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_2_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_2_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_2_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_2_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_2_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_2_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_2_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_2_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_2_io_loopExit_0_bits_control)
  );
  LoopBlockNode_3 Loop_3 ( // @[bbgemm.scala 68:22]
    .clock(Loop_3_clock),
    .reset(Loop_3_reset),
    .io_enable_ready(Loop_3_io_enable_ready),
    .io_enable_valid(Loop_3_io_enable_valid),
    .io_enable_bits_taskID(Loop_3_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_3_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_3_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_3_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_3_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_3_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_3_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_taskID(Loop_3_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_3_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_3_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_3_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_3_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_3_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_3_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_3_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_taskID(Loop_3_io_InLiveIn_3_bits_taskID),
    .io_InLiveIn_3_bits_data(Loop_3_io_InLiveIn_3_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_3_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_3_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_taskID(Loop_3_io_OutLiveIn_field3_0_bits_taskID),
    .io_OutLiveIn_field3_0_bits_data(Loop_3_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_3_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_3_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_3_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_3_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_3_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_3_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_3_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_3_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_3_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_3_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_3_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_3_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_3_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_3_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_3_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_3_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_3_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_3_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_3_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_3_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_3_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_3_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_3_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_3_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_3_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_3_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_3_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_3_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_3_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_3_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_3_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_3_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_3_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_3_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_3_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_3_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_3_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_3_io_loopExit_0_bits_control)
  );
  LoopBlockNode_4 Loop_4 ( // @[bbgemm.scala 70:22]
    .clock(Loop_4_clock),
    .reset(Loop_4_reset),
    .io_enable_ready(Loop_4_io_enable_ready),
    .io_enable_valid(Loop_4_io_enable_valid),
    .io_enable_bits_taskID(Loop_4_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_4_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_4_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_4_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_taskID(Loop_4_io_InLiveIn_0_bits_taskID),
    .io_InLiveIn_0_bits_data(Loop_4_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_4_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_4_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_taskID(Loop_4_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_4_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_4_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_4_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_4_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_4_io_InLiveIn_2_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_4_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_4_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_4_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_4_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_4_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_4_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_4_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_4_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_4_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_4_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_taskID(Loop_4_io_OutLiveIn_field0_0_bits_taskID),
    .io_OutLiveIn_field0_0_bits_data(Loop_4_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_4_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_4_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_4_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_4_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_4_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_4_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_4_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_4_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_4_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_4_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_4_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_4_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_4_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_4_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_4_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_4_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_4_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_4_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_4_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_4_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_4_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_4_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_4_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_4_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_4_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_4_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_4_io_loopExit_0_bits_control)
  );
  BasicBlockNoMaskFastNode bb_0 ( // @[bbgemm.scala 78:20]
    .clock(bb_0_clock),
    .reset(bb_0_reset),
    .io_predicateIn_0_ready(bb_0_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_0_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_0_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_0_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_0_io_Out_0_ready),
    .io_Out_0_valid(bb_0_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_0_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_0_io_Out_0_bits_control)
  );
  BasicBlockNode bb_1 ( // @[bbgemm.scala 80:20]
    .clock(bb_1_clock),
    .reset(bb_1_reset),
    .io_MaskBB_0_ready(bb_1_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_1_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_1_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_1_io_Out_0_ready),
    .io_Out_0_valid(bb_1_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_1_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_1_io_Out_1_ready),
    .io_Out_1_valid(bb_1_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_1_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_1_io_Out_1_bits_control),
    .io_Out_2_ready(bb_1_io_Out_2_ready),
    .io_Out_2_valid(bb_1_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_1_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_1_io_Out_2_bits_control),
    .io_predicateIn_0_ready(bb_1_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_1_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_1_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_1_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_1_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_1_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_1_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_1_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_1 bb_2 ( // @[bbgemm.scala 82:20]
    .clock(bb_2_clock),
    .reset(bb_2_reset),
    .io_MaskBB_0_ready(bb_2_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_2_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_2_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_2_io_Out_0_ready),
    .io_Out_0_valid(bb_2_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_2_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_2_io_Out_1_ready),
    .io_Out_1_valid(bb_2_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_2_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_2_io_Out_1_bits_control),
    .io_Out_2_ready(bb_2_io_Out_2_ready),
    .io_Out_2_valid(bb_2_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_2_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_2_io_Out_2_bits_control),
    .io_predicateIn_0_ready(bb_2_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_2_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_2_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_2_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_2_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_2_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_2_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_2_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_2 bb_3 ( // @[bbgemm.scala 84:20]
    .clock(bb_3_clock),
    .reset(bb_3_reset),
    .io_MaskBB_0_ready(bb_3_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_3_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_3_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_3_io_Out_0_ready),
    .io_Out_0_valid(bb_3_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_3_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_3_io_Out_1_ready),
    .io_Out_1_valid(bb_3_io_Out_1_valid),
    .io_Out_2_ready(bb_3_io_Out_2_ready),
    .io_Out_2_valid(bb_3_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_3_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_3_io_Out_2_bits_control),
    .io_Out_3_ready(bb_3_io_Out_3_ready),
    .io_Out_3_valid(bb_3_io_Out_3_valid),
    .io_Out_3_bits_control(bb_3_io_Out_3_bits_control),
    .io_Out_4_ready(bb_3_io_Out_4_ready),
    .io_Out_4_valid(bb_3_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_3_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_3_io_Out_4_bits_control),
    .io_predicateIn_0_ready(bb_3_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_3_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_3_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_3_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_3_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_3_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_3_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_3_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_3 bb_4 ( // @[bbgemm.scala 86:20]
    .clock(bb_4_clock),
    .reset(bb_4_reset),
    .io_MaskBB_0_ready(bb_4_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_4_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_4_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_4_io_Out_0_ready),
    .io_Out_0_valid(bb_4_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_4_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_4_io_Out_1_ready),
    .io_Out_1_valid(bb_4_io_Out_1_valid),
    .io_Out_2_ready(bb_4_io_Out_2_ready),
    .io_Out_2_valid(bb_4_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_4_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_4_io_Out_2_bits_control),
    .io_Out_3_ready(bb_4_io_Out_3_ready),
    .io_Out_3_valid(bb_4_io_Out_3_valid),
    .io_Out_3_bits_control(bb_4_io_Out_3_bits_control),
    .io_Out_4_ready(bb_4_io_Out_4_ready),
    .io_Out_4_valid(bb_4_io_Out_4_valid),
    .io_Out_4_bits_control(bb_4_io_Out_4_bits_control),
    .io_Out_5_ready(bb_4_io_Out_5_ready),
    .io_Out_5_valid(bb_4_io_Out_5_valid),
    .io_Out_5_bits_control(bb_4_io_Out_5_bits_control),
    .io_Out_6_ready(bb_4_io_Out_6_ready),
    .io_Out_6_valid(bb_4_io_Out_6_valid),
    .io_Out_6_bits_control(bb_4_io_Out_6_bits_control),
    .io_Out_7_ready(bb_4_io_Out_7_ready),
    .io_Out_7_valid(bb_4_io_Out_7_valid),
    .io_Out_7_bits_control(bb_4_io_Out_7_bits_control),
    .io_Out_8_ready(bb_4_io_Out_8_ready),
    .io_Out_8_valid(bb_4_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_4_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_4_io_Out_8_bits_control),
    .io_Out_9_ready(bb_4_io_Out_9_ready),
    .io_Out_9_valid(bb_4_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_4_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_4_io_Out_9_bits_control),
    .io_predicateIn_0_ready(bb_4_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_4_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_4_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_4_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_4_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_4_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_4_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_4_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_4 bb_5 ( // @[bbgemm.scala 88:20]
    .clock(bb_5_clock),
    .reset(bb_5_reset),
    .io_MaskBB_0_ready(bb_5_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_5_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_5_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_5_io_Out_0_ready),
    .io_Out_0_valid(bb_5_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_5_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_5_io_Out_1_ready),
    .io_Out_1_valid(bb_5_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_5_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_5_io_Out_2_ready),
    .io_Out_2_valid(bb_5_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_5_io_Out_2_bits_taskID),
    .io_Out_3_ready(bb_5_io_Out_3_ready),
    .io_Out_3_valid(bb_5_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_5_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_5_io_Out_3_bits_control),
    .io_Out_4_ready(bb_5_io_Out_4_ready),
    .io_Out_4_valid(bb_5_io_Out_4_valid),
    .io_Out_4_bits_control(bb_5_io_Out_4_bits_control),
    .io_Out_5_ready(bb_5_io_Out_5_ready),
    .io_Out_5_valid(bb_5_io_Out_5_valid),
    .io_Out_5_bits_control(bb_5_io_Out_5_bits_control),
    .io_Out_6_ready(bb_5_io_Out_6_ready),
    .io_Out_6_valid(bb_5_io_Out_6_valid),
    .io_Out_6_bits_control(bb_5_io_Out_6_bits_control),
    .io_Out_7_ready(bb_5_io_Out_7_ready),
    .io_Out_7_valid(bb_5_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_5_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_5_io_Out_7_bits_control),
    .io_Out_8_ready(bb_5_io_Out_8_ready),
    .io_Out_8_valid(bb_5_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_5_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_5_io_Out_8_bits_control),
    .io_Out_9_ready(bb_5_io_Out_9_ready),
    .io_Out_9_valid(bb_5_io_Out_9_valid),
    .io_Out_9_bits_control(bb_5_io_Out_9_bits_control),
    .io_Out_10_ready(bb_5_io_Out_10_ready),
    .io_Out_10_valid(bb_5_io_Out_10_valid),
    .io_Out_10_bits_control(bb_5_io_Out_10_bits_control),
    .io_Out_11_ready(bb_5_io_Out_11_ready),
    .io_Out_11_valid(bb_5_io_Out_11_valid),
    .io_Out_11_bits_control(bb_5_io_Out_11_bits_control),
    .io_Out_12_ready(bb_5_io_Out_12_ready),
    .io_Out_12_valid(bb_5_io_Out_12_valid),
    .io_Out_12_bits_taskID(bb_5_io_Out_12_bits_taskID),
    .io_Out_12_bits_control(bb_5_io_Out_12_bits_control),
    .io_Out_13_ready(bb_5_io_Out_13_ready),
    .io_Out_13_valid(bb_5_io_Out_13_valid),
    .io_Out_13_bits_taskID(bb_5_io_Out_13_bits_taskID),
    .io_Out_13_bits_control(bb_5_io_Out_13_bits_control),
    .io_Out_14_ready(bb_5_io_Out_14_ready),
    .io_Out_14_valid(bb_5_io_Out_14_valid),
    .io_Out_14_bits_taskID(bb_5_io_Out_14_bits_taskID),
    .io_Out_14_bits_control(bb_5_io_Out_14_bits_control),
    .io_Out_15_ready(bb_5_io_Out_15_ready),
    .io_Out_15_valid(bb_5_io_Out_15_valid),
    .io_Out_15_bits_taskID(bb_5_io_Out_15_bits_taskID),
    .io_Out_15_bits_control(bb_5_io_Out_15_bits_control),
    .io_Out_16_ready(bb_5_io_Out_16_ready),
    .io_Out_16_valid(bb_5_io_Out_16_valid),
    .io_Out_16_bits_taskID(bb_5_io_Out_16_bits_taskID),
    .io_Out_16_bits_control(bb_5_io_Out_16_bits_control),
    .io_Out_17_ready(bb_5_io_Out_17_ready),
    .io_Out_17_valid(bb_5_io_Out_17_valid),
    .io_Out_17_bits_taskID(bb_5_io_Out_17_bits_taskID),
    .io_Out_17_bits_control(bb_5_io_Out_17_bits_control),
    .io_predicateIn_0_ready(bb_5_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_5_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_5_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_5_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_5_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_5_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_5_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_5_io_predicateIn_1_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_6 ( // @[bbgemm.scala 90:20]
    .clock(bb_6_clock),
    .reset(bb_6_reset),
    .io_predicateIn_0_ready(bb_6_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_6_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_6_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_6_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_6_io_Out_0_ready),
    .io_Out_0_valid(bb_6_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_6_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_6_io_Out_1_ready),
    .io_Out_1_valid(bb_6_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_6_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_6_io_Out_2_ready),
    .io_Out_2_valid(bb_6_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_6_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_6_io_Out_2_bits_control),
    .io_Out_3_ready(bb_6_io_Out_3_ready),
    .io_Out_3_valid(bb_6_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_6_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_6_io_Out_3_bits_control),
    .io_Out_4_ready(bb_6_io_Out_4_ready),
    .io_Out_4_valid(bb_6_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_6_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_6_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_7 ( // @[bbgemm.scala 92:20]
    .clock(bb_7_clock),
    .reset(bb_7_reset),
    .io_predicateIn_0_ready(bb_7_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_7_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_7_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_7_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_7_io_Out_0_ready),
    .io_Out_0_valid(bb_7_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_7_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_7_io_Out_1_ready),
    .io_Out_1_valid(bb_7_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_7_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_7_io_Out_2_ready),
    .io_Out_2_valid(bb_7_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_7_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_7_io_Out_2_bits_control),
    .io_Out_3_ready(bb_7_io_Out_3_ready),
    .io_Out_3_valid(bb_7_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_7_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_7_io_Out_3_bits_control),
    .io_Out_4_ready(bb_7_io_Out_4_ready),
    .io_Out_4_valid(bb_7_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_7_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_7_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_8 ( // @[bbgemm.scala 94:20]
    .clock(bb_8_clock),
    .reset(bb_8_reset),
    .io_predicateIn_0_ready(bb_8_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_8_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_8_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_8_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_8_io_Out_0_ready),
    .io_Out_0_valid(bb_8_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_8_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_8_io_Out_1_ready),
    .io_Out_1_valid(bb_8_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_8_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_8_io_Out_2_ready),
    .io_Out_2_valid(bb_8_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_8_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_8_io_Out_2_bits_control),
    .io_Out_3_ready(bb_8_io_Out_3_ready),
    .io_Out_3_valid(bb_8_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_8_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_8_io_Out_3_bits_control),
    .io_Out_4_ready(bb_8_io_Out_4_ready),
    .io_Out_4_valid(bb_8_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_8_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_8_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_9 ( // @[bbgemm.scala 96:20]
    .clock(bb_9_clock),
    .reset(bb_9_reset),
    .io_predicateIn_0_ready(bb_9_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_9_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_9_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_9_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_9_io_Out_0_ready),
    .io_Out_0_valid(bb_9_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_9_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_9_io_Out_1_ready),
    .io_Out_1_valid(bb_9_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_9_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_9_io_Out_2_ready),
    .io_Out_2_valid(bb_9_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_9_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_9_io_Out_2_bits_control),
    .io_Out_3_ready(bb_9_io_Out_3_ready),
    .io_Out_3_valid(bb_9_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_9_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_9_io_Out_3_bits_control),
    .io_Out_4_ready(bb_9_io_Out_4_ready),
    .io_Out_4_valid(bb_9_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_9_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_9_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode bb_10 ( // @[bbgemm.scala 98:21]
    .clock(bb_10_clock),
    .reset(bb_10_reset),
    .io_predicateIn_0_ready(bb_10_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_10_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_10_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_10_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_10_io_Out_0_ready),
    .io_Out_0_valid(bb_10_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_10_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_10_io_Out_0_bits_control)
  );
  UBranchNode br_0 ( // @[bbgemm.scala 107:20]
    .clock(br_0_clock),
    .reset(br_0_reset),
    .io_enable_ready(br_0_io_enable_ready),
    .io_enable_valid(br_0_io_enable_valid),
    .io_enable_bits_taskID(br_0_io_enable_bits_taskID),
    .io_enable_bits_control(br_0_io_enable_bits_control),
    .io_Out_0_ready(br_0_io_Out_0_ready),
    .io_Out_0_valid(br_0_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_0_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_0_io_Out_0_bits_control)
  );
  PhiFastNode phi1 ( // @[bbgemm.scala 110:20]
    .clock(phi1_clock),
    .reset(phi1_reset),
    .io_enable_ready(phi1_io_enable_ready),
    .io_enable_valid(phi1_io_enable_valid),
    .io_enable_bits_taskID(phi1_io_enable_bits_taskID),
    .io_enable_bits_control(phi1_io_enable_bits_control),
    .io_InData_0_ready(phi1_io_InData_0_ready),
    .io_InData_0_valid(phi1_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi1_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi1_io_InData_1_ready),
    .io_InData_1_valid(phi1_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi1_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi1_io_InData_1_bits_data),
    .io_Mask_ready(phi1_io_Mask_ready),
    .io_Mask_valid(phi1_io_Mask_valid),
    .io_Mask_bits(phi1_io_Mask_bits),
    .io_Out_0_ready(phi1_io_Out_0_ready),
    .io_Out_0_valid(phi1_io_Out_0_valid),
    .io_Out_0_bits_data(phi1_io_Out_0_bits_data),
    .io_Out_1_ready(phi1_io_Out_1_ready),
    .io_Out_1_valid(phi1_io_Out_1_valid),
    .io_Out_1_bits_taskID(phi1_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(phi1_io_Out_1_bits_data)
  );
  UBranchNode_1 br_2 ( // @[bbgemm.scala 113:20]
    .clock(br_2_clock),
    .reset(br_2_reset),
    .io_enable_ready(br_2_io_enable_ready),
    .io_enable_valid(br_2_io_enable_valid),
    .io_enable_bits_taskID(br_2_io_enable_bits_taskID),
    .io_enable_bits_control(br_2_io_enable_bits_control),
    .io_Out_0_ready(br_2_io_Out_0_ready),
    .io_Out_0_valid(br_2_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_2_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_2_io_Out_0_bits_control)
  );
  PhiFastNode phi3 ( // @[bbgemm.scala 116:20]
    .clock(phi3_clock),
    .reset(phi3_reset),
    .io_enable_ready(phi3_io_enable_ready),
    .io_enable_valid(phi3_io_enable_valid),
    .io_enable_bits_taskID(phi3_io_enable_bits_taskID),
    .io_enable_bits_control(phi3_io_enable_bits_control),
    .io_InData_0_ready(phi3_io_InData_0_ready),
    .io_InData_0_valid(phi3_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi3_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi3_io_InData_1_ready),
    .io_InData_1_valid(phi3_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi3_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi3_io_InData_1_bits_data),
    .io_Mask_ready(phi3_io_Mask_ready),
    .io_Mask_valid(phi3_io_Mask_valid),
    .io_Mask_bits(phi3_io_Mask_bits),
    .io_Out_0_ready(phi3_io_Out_0_ready),
    .io_Out_0_valid(phi3_io_Out_0_valid),
    .io_Out_0_bits_data(phi3_io_Out_0_bits_data),
    .io_Out_1_ready(phi3_io_Out_1_ready),
    .io_Out_1_valid(phi3_io_Out_1_valid),
    .io_Out_1_bits_taskID(phi3_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(phi3_io_Out_1_bits_data)
  );
  UBranchNode_2 br_4 ( // @[bbgemm.scala 119:20]
    .clock(br_4_clock),
    .reset(br_4_reset),
    .io_enable_ready(br_4_io_enable_ready),
    .io_enable_valid(br_4_io_enable_valid),
    .io_enable_bits_taskID(br_4_io_enable_bits_taskID),
    .io_enable_bits_control(br_4_io_enable_bits_control),
    .io_Out_0_ready(br_4_io_Out_0_ready),
    .io_Out_0_valid(br_4_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_4_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_4_io_Out_0_bits_control)
  );
  PhiFastNode_2 phi5 ( // @[bbgemm.scala 122:20]
    .clock(phi5_clock),
    .reset(phi5_reset),
    .io_enable_ready(phi5_io_enable_ready),
    .io_enable_valid(phi5_io_enable_valid),
    .io_enable_bits_taskID(phi5_io_enable_bits_taskID),
    .io_enable_bits_control(phi5_io_enable_bits_control),
    .io_InData_0_ready(phi5_io_InData_0_ready),
    .io_InData_0_valid(phi5_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi5_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi5_io_InData_1_ready),
    .io_InData_1_valid(phi5_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi5_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi5_io_InData_1_bits_data),
    .io_Mask_ready(phi5_io_Mask_ready),
    .io_Mask_valid(phi5_io_Mask_valid),
    .io_Mask_bits(phi5_io_Mask_bits),
    .io_Out_0_ready(phi5_io_Out_0_ready),
    .io_Out_0_valid(phi5_io_Out_0_valid),
    .io_Out_0_bits_data(phi5_io_Out_0_bits_data),
    .io_Out_1_ready(phi5_io_Out_1_ready),
    .io_Out_1_valid(phi5_io_Out_1_valid),
    .io_Out_1_bits_taskID(phi5_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(phi5_io_Out_1_bits_data)
  );
  ComputeNode binaryOp_6 ( // @[bbgemm.scala 125:26]
    .clock(binaryOp_6_clock),
    .reset(binaryOp_6_reset),
    .io_enable_ready(binaryOp_6_io_enable_ready),
    .io_enable_valid(binaryOp_6_io_enable_valid),
    .io_enable_bits_control(binaryOp_6_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_6_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_6_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_6_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_6_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_6_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_6_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_6_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_6_io_RightIO_valid)
  );
  UBranchNode_3 br_7 ( // @[bbgemm.scala 128:20]
    .clock(br_7_clock),
    .reset(br_7_reset),
    .io_enable_ready(br_7_io_enable_ready),
    .io_enable_valid(br_7_io_enable_valid),
    .io_enable_bits_taskID(br_7_io_enable_bits_taskID),
    .io_enable_bits_control(br_7_io_enable_bits_control),
    .io_Out_0_ready(br_7_io_Out_0_ready),
    .io_Out_0_valid(br_7_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_7_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_7_io_Out_0_bits_control)
  );
  PhiFastNode_3 phi8 ( // @[bbgemm.scala 131:20]
    .clock(phi8_clock),
    .reset(phi8_reset),
    .io_enable_ready(phi8_io_enable_ready),
    .io_enable_valid(phi8_io_enable_valid),
    .io_enable_bits_taskID(phi8_io_enable_bits_taskID),
    .io_enable_bits_control(phi8_io_enable_bits_control),
    .io_InData_0_ready(phi8_io_InData_0_ready),
    .io_InData_0_valid(phi8_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi8_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi8_io_InData_1_ready),
    .io_InData_1_valid(phi8_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi8_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi8_io_InData_1_bits_data),
    .io_Mask_ready(phi8_io_Mask_ready),
    .io_Mask_valid(phi8_io_Mask_valid),
    .io_Mask_bits(phi8_io_Mask_bits),
    .io_Out_0_ready(phi8_io_Out_0_ready),
    .io_Out_0_valid(phi8_io_Out_0_valid),
    .io_Out_0_bits_data(phi8_io_Out_0_bits_data),
    .io_Out_1_ready(phi8_io_Out_1_ready),
    .io_Out_1_valid(phi8_io_Out_1_valid),
    .io_Out_1_bits_data(phi8_io_Out_1_bits_data),
    .io_Out_2_ready(phi8_io_Out_2_ready),
    .io_Out_2_valid(phi8_io_Out_2_valid),
    .io_Out_2_bits_taskID(phi8_io_Out_2_bits_taskID),
    .io_Out_2_bits_data(phi8_io_Out_2_bits_data)
  );
  ComputeNode_1 binaryOp_9 ( // @[bbgemm.scala 134:26]
    .clock(binaryOp_9_clock),
    .reset(binaryOp_9_reset),
    .io_enable_ready(binaryOp_9_io_enable_ready),
    .io_enable_valid(binaryOp_9_io_enable_valid),
    .io_enable_bits_control(binaryOp_9_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_9_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_9_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_9_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_9_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_9_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_9_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_9_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_9_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_9_io_RightIO_bits_data)
  );
  ComputeNode_2 binaryOp_10 ( // @[bbgemm.scala 137:27]
    .clock(binaryOp_10_clock),
    .reset(binaryOp_10_reset),
    .io_enable_ready(binaryOp_10_io_enable_ready),
    .io_enable_valid(binaryOp_10_io_enable_valid),
    .io_enable_bits_control(binaryOp_10_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_10_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_10_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_10_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_10_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_10_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_10_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_10_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_10_io_RightIO_valid)
  );
  ComputeNode_3 binaryOp_11 ( // @[bbgemm.scala 140:27]
    .clock(binaryOp_11_clock),
    .reset(binaryOp_11_reset),
    .io_enable_ready(binaryOp_11_io_enable_ready),
    .io_enable_valid(binaryOp_11_io_enable_valid),
    .io_enable_bits_control(binaryOp_11_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_11_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_11_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_11_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_11_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_11_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_11_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_11_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_11_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_11_io_RightIO_bits_data)
  );
  ComputeNode_4 binaryOp_12 ( // @[bbgemm.scala 143:27]
    .clock(binaryOp_12_clock),
    .reset(binaryOp_12_reset),
    .io_enable_ready(binaryOp_12_io_enable_ready),
    .io_enable_valid(binaryOp_12_io_enable_valid),
    .io_enable_bits_control(binaryOp_12_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_12_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_12_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_12_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_12_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_12_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_12_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_12_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_12_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_12_io_RightIO_bits_data)
  );
  GepNode Gep_13 ( // @[bbgemm.scala 146:22]
    .clock(Gep_13_clock),
    .reset(Gep_13_reset),
    .io_enable_ready(Gep_13_io_enable_ready),
    .io_enable_valid(Gep_13_io_enable_valid),
    .io_enable_bits_control(Gep_13_io_enable_bits_control),
    .io_Out_0_ready(Gep_13_io_Out_0_ready),
    .io_Out_0_valid(Gep_13_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_13_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_13_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_13_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_13_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_13_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_13_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_13_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_13_io_idx_0_ready),
    .io_idx_0_valid(Gep_13_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_13_io_idx_0_bits_data)
  );
  UnTypLoad ld_14 ( // @[bbgemm.scala 149:21]
    .clock(ld_14_clock),
    .reset(ld_14_reset),
    .io_enable_ready(ld_14_io_enable_ready),
    .io_enable_valid(ld_14_io_enable_valid),
    .io_enable_bits_taskID(ld_14_io_enable_bits_taskID),
    .io_enable_bits_control(ld_14_io_enable_bits_control),
    .io_Out_0_ready(ld_14_io_Out_0_ready),
    .io_Out_0_valid(ld_14_io_Out_0_valid),
    .io_Out_0_bits_taskID(ld_14_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(ld_14_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_14_io_GepAddr_ready),
    .io_GepAddr_valid(ld_14_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_14_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_14_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_14_io_GepAddr_bits_data),
    .io_memReq_ready(ld_14_io_memReq_ready),
    .io_memReq_valid(ld_14_io_memReq_valid),
    .io_memReq_bits_address(ld_14_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_14_io_memReq_bits_taskID),
    .io_memResp_valid(ld_14_io_memResp_valid),
    .io_memResp_data(ld_14_io_memResp_data)
  );
  UBranchNode_4 br_15 ( // @[bbgemm.scala 152:21]
    .clock(br_15_clock),
    .reset(br_15_reset),
    .io_enable_ready(br_15_io_enable_ready),
    .io_enable_valid(br_15_io_enable_valid),
    .io_enable_bits_taskID(br_15_io_enable_bits_taskID),
    .io_enable_bits_control(br_15_io_enable_bits_control),
    .io_Out_0_ready(br_15_io_Out_0_ready),
    .io_Out_0_valid(br_15_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_15_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_15_io_Out_0_bits_control)
  );
  PhiFastNode_3 phi16 ( // @[bbgemm.scala 155:21]
    .clock(phi16_clock),
    .reset(phi16_reset),
    .io_enable_ready(phi16_io_enable_ready),
    .io_enable_valid(phi16_io_enable_valid),
    .io_enable_bits_taskID(phi16_io_enable_bits_taskID),
    .io_enable_bits_control(phi16_io_enable_bits_control),
    .io_InData_0_ready(phi16_io_InData_0_ready),
    .io_InData_0_valid(phi16_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi16_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi16_io_InData_1_ready),
    .io_InData_1_valid(phi16_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi16_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi16_io_InData_1_bits_data),
    .io_Mask_ready(phi16_io_Mask_ready),
    .io_Mask_valid(phi16_io_Mask_valid),
    .io_Mask_bits(phi16_io_Mask_bits),
    .io_Out_0_ready(phi16_io_Out_0_ready),
    .io_Out_0_valid(phi16_io_Out_0_valid),
    .io_Out_0_bits_data(phi16_io_Out_0_bits_data),
    .io_Out_1_ready(phi16_io_Out_1_ready),
    .io_Out_1_valid(phi16_io_Out_1_valid),
    .io_Out_1_bits_data(phi16_io_Out_1_bits_data),
    .io_Out_2_ready(phi16_io_Out_2_ready),
    .io_Out_2_valid(phi16_io_Out_2_valid),
    .io_Out_2_bits_taskID(phi16_io_Out_2_bits_taskID),
    .io_Out_2_bits_data(phi16_io_Out_2_bits_data)
  );
  ComputeNode_5 binaryOp_17 ( // @[bbgemm.scala 158:27]
    .clock(binaryOp_17_clock),
    .reset(binaryOp_17_reset),
    .io_enable_ready(binaryOp_17_io_enable_ready),
    .io_enable_valid(binaryOp_17_io_enable_valid),
    .io_enable_bits_control(binaryOp_17_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_17_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_17_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_17_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_17_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_17_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_17_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_17_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_17_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_17_io_RightIO_bits_data)
  );
  ComputeNode_6 binaryOp_18 ( // @[bbgemm.scala 161:27]
    .clock(binaryOp_18_clock),
    .reset(binaryOp_18_reset),
    .io_enable_ready(binaryOp_18_io_enable_ready),
    .io_enable_valid(binaryOp_18_io_enable_valid),
    .io_enable_bits_control(binaryOp_18_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_18_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_18_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_18_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_18_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_18_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_18_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_18_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_18_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_18_io_RightIO_bits_data)
  );
  GepNode_1 Gep_19 ( // @[bbgemm.scala 164:22]
    .clock(Gep_19_clock),
    .reset(Gep_19_reset),
    .io_enable_ready(Gep_19_io_enable_ready),
    .io_enable_valid(Gep_19_io_enable_valid),
    .io_enable_bits_control(Gep_19_io_enable_bits_control),
    .io_Out_0_ready(Gep_19_io_Out_0_ready),
    .io_Out_0_valid(Gep_19_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_19_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_19_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_19_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_19_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_19_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_19_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_19_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_19_io_idx_0_ready),
    .io_idx_0_valid(Gep_19_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_19_io_idx_0_bits_data)
  );
  UnTypLoad_1 ld_20 ( // @[bbgemm.scala 167:21]
    .clock(ld_20_clock),
    .reset(ld_20_reset),
    .io_enable_ready(ld_20_io_enable_ready),
    .io_enable_valid(ld_20_io_enable_valid),
    .io_enable_bits_taskID(ld_20_io_enable_bits_taskID),
    .io_enable_bits_control(ld_20_io_enable_bits_control),
    .io_Out_0_ready(ld_20_io_Out_0_ready),
    .io_Out_0_valid(ld_20_io_Out_0_valid),
    .io_Out_0_bits_taskID(ld_20_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(ld_20_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_20_io_GepAddr_ready),
    .io_GepAddr_valid(ld_20_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_20_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_20_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_20_io_GepAddr_bits_data),
    .io_memReq_ready(ld_20_io_memReq_ready),
    .io_memReq_valid(ld_20_io_memReq_valid),
    .io_memReq_bits_address(ld_20_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_20_io_memReq_bits_taskID),
    .io_memResp_valid(ld_20_io_memResp_valid),
    .io_memResp_data(ld_20_io_memResp_data)
  );
  FPCustomMultiplierNode FP_21 ( // @[bbgemm.scala 171:21]
    .clock(FP_21_clock),
    .reset(FP_21_reset),
    .io_enable_ready(FP_21_io_enable_ready),
    .io_enable_valid(FP_21_io_enable_valid),
    .io_enable_bits_taskID(FP_21_io_enable_bits_taskID),
    .io_enable_bits_control(FP_21_io_enable_bits_control),
    .io_Out_0_ready(FP_21_io_Out_0_ready),
    .io_Out_0_valid(FP_21_io_Out_0_valid),
    .io_Out_0_bits_taskID(FP_21_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(FP_21_io_Out_0_bits_data),
    .io_LeftIO_ready(FP_21_io_LeftIO_ready),
    .io_LeftIO_valid(FP_21_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(FP_21_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(FP_21_io_LeftIO_bits_data),
    .io_RightIO_ready(FP_21_io_RightIO_ready),
    .io_RightIO_valid(FP_21_io_RightIO_valid),
    .io_RightIO_bits_taskID(FP_21_io_RightIO_bits_taskID),
    .io_RightIO_bits_data(FP_21_io_RightIO_bits_data)
  );
  ComputeNode_7 binaryOp_22 ( // @[bbgemm.scala 174:27]
    .clock(binaryOp_22_clock),
    .reset(binaryOp_22_reset),
    .io_enable_ready(binaryOp_22_io_enable_ready),
    .io_enable_valid(binaryOp_22_io_enable_valid),
    .io_enable_bits_control(binaryOp_22_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_22_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_22_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_22_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_22_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_22_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_22_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_22_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_22_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_22_io_RightIO_bits_data)
  );
  ComputeNode_8 binaryOp_23 ( // @[bbgemm.scala 177:27]
    .clock(binaryOp_23_clock),
    .reset(binaryOp_23_reset),
    .io_enable_ready(binaryOp_23_io_enable_ready),
    .io_enable_valid(binaryOp_23_io_enable_valid),
    .io_enable_bits_control(binaryOp_23_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_23_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_23_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_23_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_23_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_23_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_23_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_23_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_23_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_23_io_RightIO_bits_data)
  );
  GepNode_2 Gep_24 ( // @[bbgemm.scala 180:22]
    .clock(Gep_24_clock),
    .reset(Gep_24_reset),
    .io_enable_ready(Gep_24_io_enable_ready),
    .io_enable_valid(Gep_24_io_enable_valid),
    .io_enable_bits_control(Gep_24_io_enable_bits_control),
    .io_Out_0_ready(Gep_24_io_Out_0_ready),
    .io_Out_0_valid(Gep_24_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_24_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_24_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_24_io_Out_0_bits_data),
    .io_Out_1_ready(Gep_24_io_Out_1_ready),
    .io_Out_1_valid(Gep_24_io_Out_1_valid),
    .io_Out_1_bits_taskID(Gep_24_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(Gep_24_io_Out_1_bits_data),
    .io_baseAddress_ready(Gep_24_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_24_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_24_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_24_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_24_io_idx_0_ready),
    .io_idx_0_valid(Gep_24_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_24_io_idx_0_bits_data)
  );
  UnTypLoad_2 ld_25 ( // @[bbgemm.scala 183:21]
    .clock(ld_25_clock),
    .reset(ld_25_reset),
    .io_enable_ready(ld_25_io_enable_ready),
    .io_enable_valid(ld_25_io_enable_valid),
    .io_enable_bits_taskID(ld_25_io_enable_bits_taskID),
    .io_enable_bits_control(ld_25_io_enable_bits_control),
    .io_Out_0_ready(ld_25_io_Out_0_ready),
    .io_Out_0_valid(ld_25_io_Out_0_valid),
    .io_Out_0_bits_taskID(ld_25_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(ld_25_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_25_io_GepAddr_ready),
    .io_GepAddr_valid(ld_25_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_25_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_25_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_25_io_GepAddr_bits_data),
    .io_memReq_ready(ld_25_io_memReq_ready),
    .io_memReq_valid(ld_25_io_memReq_valid),
    .io_memReq_bits_address(ld_25_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_25_io_memReq_bits_taskID),
    .io_memResp_valid(ld_25_io_memResp_valid),
    .io_memResp_data(ld_25_io_memResp_data)
  );
  FPCustomAdderNode FP_26 ( // @[bbgemm.scala 187:21]
    .clock(FP_26_clock),
    .reset(FP_26_reset),
    .io_enable_ready(FP_26_io_enable_ready),
    .io_enable_valid(FP_26_io_enable_valid),
    .io_enable_bits_taskID(FP_26_io_enable_bits_taskID),
    .io_enable_bits_control(FP_26_io_enable_bits_control),
    .io_Out_0_ready(FP_26_io_Out_0_ready),
    .io_Out_0_valid(FP_26_io_Out_0_valid),
    .io_Out_0_bits_taskID(FP_26_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(FP_26_io_Out_0_bits_data),
    .io_LeftIO_ready(FP_26_io_LeftIO_ready),
    .io_LeftIO_valid(FP_26_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(FP_26_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(FP_26_io_LeftIO_bits_data),
    .io_RightIO_ready(FP_26_io_RightIO_ready),
    .io_RightIO_valid(FP_26_io_RightIO_valid),
    .io_RightIO_bits_taskID(FP_26_io_RightIO_bits_taskID),
    .io_RightIO_bits_data(FP_26_io_RightIO_bits_data)
  );
  UnTypStore st_27 ( // @[bbgemm.scala 190:21]
    .clock(st_27_clock),
    .reset(st_27_reset),
    .io_enable_ready(st_27_io_enable_ready),
    .io_enable_valid(st_27_io_enable_valid),
    .io_enable_bits_taskID(st_27_io_enable_bits_taskID),
    .io_enable_bits_control(st_27_io_enable_bits_control),
    .io_GepAddr_ready(st_27_io_GepAddr_ready),
    .io_GepAddr_valid(st_27_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_27_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_27_io_GepAddr_bits_data),
    .io_inData_ready(st_27_io_inData_ready),
    .io_inData_valid(st_27_io_inData_valid),
    .io_inData_bits_taskID(st_27_io_inData_bits_taskID),
    .io_inData_bits_data(st_27_io_inData_bits_data),
    .io_memReq_ready(st_27_io_memReq_ready),
    .io_memReq_valid(st_27_io_memReq_valid),
    .io_memReq_bits_address(st_27_io_memReq_bits_address),
    .io_memReq_bits_data(st_27_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_27_io_memReq_bits_taskID),
    .io_memResp_valid(st_27_io_memResp_valid)
  );
  ComputeNode_9 binaryOp_28 ( // @[bbgemm.scala 193:27]
    .clock(binaryOp_28_clock),
    .reset(binaryOp_28_reset),
    .io_enable_ready(binaryOp_28_io_enable_ready),
    .io_enable_valid(binaryOp_28_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_28_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_28_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_28_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_28_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_28_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_28_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_28_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_28_io_Out_1_valid),
    .io_Out_1_bits_taskID(binaryOp_28_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(binaryOp_28_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_28_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_28_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(binaryOp_28_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(binaryOp_28_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_28_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_28_io_RightIO_valid),
    .io_RightIO_bits_taskID(binaryOp_28_io_RightIO_bits_taskID)
  );
  IcmpNode icmp_29 ( // @[bbgemm.scala 196:23]
    .clock(icmp_29_clock),
    .reset(icmp_29_reset),
    .io_enable_ready(icmp_29_io_enable_ready),
    .io_enable_valid(icmp_29_io_enable_valid),
    .io_enable_bits_taskID(icmp_29_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_29_io_enable_bits_control),
    .io_Out_0_ready(icmp_29_io_Out_0_ready),
    .io_Out_0_valid(icmp_29_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_29_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_29_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_29_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_29_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(icmp_29_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(icmp_29_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_29_io_RightIO_ready),
    .io_RightIO_valid(icmp_29_io_RightIO_valid),
    .io_RightIO_bits_taskID(icmp_29_io_RightIO_bits_taskID)
  );
  CBranchNodeVariable br_30 ( // @[bbgemm.scala 199:21]
    .clock(br_30_clock),
    .reset(br_30_reset),
    .io_enable_ready(br_30_io_enable_ready),
    .io_enable_valid(br_30_io_enable_valid),
    .io_enable_bits_taskID(br_30_io_enable_bits_taskID),
    .io_enable_bits_control(br_30_io_enable_bits_control),
    .io_CmpIO_ready(br_30_io_CmpIO_ready),
    .io_CmpIO_valid(br_30_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_30_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_30_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_30_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_30_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_30_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_30_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_30_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_30_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_30_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_30_io_FalseOutput_0_bits_control)
  );
  ComputeNode_10 binaryOp_31 ( // @[bbgemm.scala 202:27]
    .clock(binaryOp_31_clock),
    .reset(binaryOp_31_reset),
    .io_enable_ready(binaryOp_31_io_enable_ready),
    .io_enable_valid(binaryOp_31_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_31_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_31_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_31_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_31_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_31_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_31_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_31_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_31_io_Out_1_valid),
    .io_Out_1_bits_taskID(binaryOp_31_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(binaryOp_31_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_31_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_31_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(binaryOp_31_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(binaryOp_31_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_31_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_31_io_RightIO_valid),
    .io_RightIO_bits_taskID(binaryOp_31_io_RightIO_bits_taskID)
  );
  IcmpNode_1 icmp_32 ( // @[bbgemm.scala 205:23]
    .clock(icmp_32_clock),
    .reset(icmp_32_reset),
    .io_enable_ready(icmp_32_io_enable_ready),
    .io_enable_valid(icmp_32_io_enable_valid),
    .io_enable_bits_taskID(icmp_32_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_32_io_enable_bits_control),
    .io_Out_0_ready(icmp_32_io_Out_0_ready),
    .io_Out_0_valid(icmp_32_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_32_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_32_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_32_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_32_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(icmp_32_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(icmp_32_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_32_io_RightIO_ready),
    .io_RightIO_valid(icmp_32_io_RightIO_valid),
    .io_RightIO_bits_taskID(icmp_32_io_RightIO_bits_taskID)
  );
  CBranchNodeVariable br_33 ( // @[bbgemm.scala 208:21]
    .clock(br_33_clock),
    .reset(br_33_reset),
    .io_enable_ready(br_33_io_enable_ready),
    .io_enable_valid(br_33_io_enable_valid),
    .io_enable_bits_taskID(br_33_io_enable_bits_taskID),
    .io_enable_bits_control(br_33_io_enable_bits_control),
    .io_CmpIO_ready(br_33_io_CmpIO_ready),
    .io_CmpIO_valid(br_33_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_33_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_33_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_33_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_33_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_33_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_33_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_33_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_33_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_33_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_33_io_FalseOutput_0_bits_control)
  );
  ComputeNode_11 binaryOp_34 ( // @[bbgemm.scala 211:27]
    .clock(binaryOp_34_clock),
    .reset(binaryOp_34_reset),
    .io_enable_ready(binaryOp_34_io_enable_ready),
    .io_enable_valid(binaryOp_34_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_34_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_34_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_34_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_34_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_34_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_34_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_34_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_34_io_Out_1_valid),
    .io_Out_1_bits_taskID(binaryOp_34_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(binaryOp_34_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_34_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_34_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(binaryOp_34_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(binaryOp_34_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_34_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_34_io_RightIO_valid),
    .io_RightIO_bits_taskID(binaryOp_34_io_RightIO_bits_taskID)
  );
  IcmpNode_2 icmp_35 ( // @[bbgemm.scala 214:23]
    .clock(icmp_35_clock),
    .reset(icmp_35_reset),
    .io_enable_ready(icmp_35_io_enable_ready),
    .io_enable_valid(icmp_35_io_enable_valid),
    .io_enable_bits_taskID(icmp_35_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_35_io_enable_bits_control),
    .io_Out_0_ready(icmp_35_io_Out_0_ready),
    .io_Out_0_valid(icmp_35_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_35_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_35_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_35_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_35_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(icmp_35_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(icmp_35_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_35_io_RightIO_ready),
    .io_RightIO_valid(icmp_35_io_RightIO_valid),
    .io_RightIO_bits_taskID(icmp_35_io_RightIO_bits_taskID)
  );
  CBranchNodeVariable br_36 ( // @[bbgemm.scala 217:21]
    .clock(br_36_clock),
    .reset(br_36_reset),
    .io_enable_ready(br_36_io_enable_ready),
    .io_enable_valid(br_36_io_enable_valid),
    .io_enable_bits_taskID(br_36_io_enable_bits_taskID),
    .io_enable_bits_control(br_36_io_enable_bits_control),
    .io_CmpIO_ready(br_36_io_CmpIO_ready),
    .io_CmpIO_valid(br_36_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_36_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_36_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_36_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_36_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_36_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_36_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_36_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_36_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_36_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_36_io_FalseOutput_0_bits_control)
  );
  ComputeNode_12 binaryOp_37 ( // @[bbgemm.scala 220:27]
    .clock(binaryOp_37_clock),
    .reset(binaryOp_37_reset),
    .io_enable_ready(binaryOp_37_io_enable_ready),
    .io_enable_valid(binaryOp_37_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_37_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_37_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_37_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_37_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_37_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_37_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_37_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_37_io_Out_1_valid),
    .io_Out_1_bits_taskID(binaryOp_37_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(binaryOp_37_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_37_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_37_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(binaryOp_37_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(binaryOp_37_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_37_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_37_io_RightIO_valid),
    .io_RightIO_bits_taskID(binaryOp_37_io_RightIO_bits_taskID)
  );
  IcmpNode_3 icmp_38 ( // @[bbgemm.scala 223:23]
    .clock(icmp_38_clock),
    .reset(icmp_38_reset),
    .io_enable_ready(icmp_38_io_enable_ready),
    .io_enable_valid(icmp_38_io_enable_valid),
    .io_enable_bits_taskID(icmp_38_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_38_io_enable_bits_control),
    .io_Out_0_ready(icmp_38_io_Out_0_ready),
    .io_Out_0_valid(icmp_38_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_38_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_38_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_38_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_38_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(icmp_38_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(icmp_38_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_38_io_RightIO_ready),
    .io_RightIO_valid(icmp_38_io_RightIO_valid),
    .io_RightIO_bits_taskID(icmp_38_io_RightIO_bits_taskID)
  );
  CBranchNodeVariable br_39 ( // @[bbgemm.scala 226:21]
    .clock(br_39_clock),
    .reset(br_39_reset),
    .io_enable_ready(br_39_io_enable_ready),
    .io_enable_valid(br_39_io_enable_valid),
    .io_enable_bits_taskID(br_39_io_enable_bits_taskID),
    .io_enable_bits_control(br_39_io_enable_bits_control),
    .io_CmpIO_ready(br_39_io_CmpIO_ready),
    .io_CmpIO_valid(br_39_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_39_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_39_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_39_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_39_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_39_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_39_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_39_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_39_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_39_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_39_io_FalseOutput_0_bits_control)
  );
  ComputeNode_13 binaryOp_40 ( // @[bbgemm.scala 229:27]
    .clock(binaryOp_40_clock),
    .reset(binaryOp_40_reset),
    .io_enable_ready(binaryOp_40_io_enable_ready),
    .io_enable_valid(binaryOp_40_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_40_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_40_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_40_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_40_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_40_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_40_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_40_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_40_io_Out_1_valid),
    .io_Out_1_bits_taskID(binaryOp_40_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(binaryOp_40_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_40_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_40_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(binaryOp_40_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(binaryOp_40_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_40_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_40_io_RightIO_valid),
    .io_RightIO_bits_taskID(binaryOp_40_io_RightIO_bits_taskID)
  );
  IcmpNode_4 icmp_41 ( // @[bbgemm.scala 232:23]
    .clock(icmp_41_clock),
    .reset(icmp_41_reset),
    .io_enable_ready(icmp_41_io_enable_ready),
    .io_enable_valid(icmp_41_io_enable_valid),
    .io_enable_bits_taskID(icmp_41_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_41_io_enable_bits_control),
    .io_Out_0_ready(icmp_41_io_Out_0_ready),
    .io_Out_0_valid(icmp_41_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_41_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_41_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_41_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_41_io_LeftIO_valid),
    .io_LeftIO_bits_taskID(icmp_41_io_LeftIO_bits_taskID),
    .io_LeftIO_bits_data(icmp_41_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_41_io_RightIO_ready),
    .io_RightIO_valid(icmp_41_io_RightIO_valid),
    .io_RightIO_bits_taskID(icmp_41_io_RightIO_bits_taskID)
  );
  CBranchNodeVariable br_42 ( // @[bbgemm.scala 235:21]
    .clock(br_42_clock),
    .reset(br_42_reset),
    .io_enable_ready(br_42_io_enable_ready),
    .io_enable_valid(br_42_io_enable_valid),
    .io_enable_bits_taskID(br_42_io_enable_bits_taskID),
    .io_enable_bits_control(br_42_io_enable_bits_control),
    .io_CmpIO_ready(br_42_io_CmpIO_ready),
    .io_CmpIO_valid(br_42_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_42_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_42_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_42_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_42_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_42_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_42_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_42_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_42_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_42_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_42_io_FalseOutput_0_bits_control)
  );
  RetNode2 ret_43 ( // @[bbgemm.scala 238:22]
    .clock(ret_43_clock),
    .reset(ret_43_reset),
    .io_In_enable_ready(ret_43_io_In_enable_ready),
    .io_In_enable_valid(ret_43_io_In_enable_valid),
    .io_In_enable_bits_taskID(ret_43_io_In_enable_bits_taskID),
    .io_In_enable_bits_control(ret_43_io_In_enable_bits_control),
    .io_Out_ready(ret_43_io_Out_ready),
    .io_Out_valid(ret_43_io_Out_valid),
    .io_Out_bits_enable_taskID(ret_43_io_Out_bits_enable_taskID),
    .io_Out_bits_enable_control(ret_43_io_Out_bits_enable_control)
  );
  ConstFastNode const0 ( // @[bbgemm.scala 247:22]
    .clock(const0_clock),
    .reset(const0_reset),
    .io_enable_ready(const0_io_enable_ready),
    .io_enable_valid(const0_io_enable_valid),
    .io_enable_bits_taskID(const0_io_enable_bits_taskID),
    .io_Out_ready(const0_io_Out_ready),
    .io_Out_valid(const0_io_Out_valid),
    .io_Out_bits_taskID(const0_io_Out_bits_taskID)
  );
  ConstFastNode const1 ( // @[bbgemm.scala 250:22]
    .clock(const1_clock),
    .reset(const1_reset),
    .io_enable_ready(const1_io_enable_ready),
    .io_enable_valid(const1_io_enable_valid),
    .io_enable_bits_taskID(const1_io_enable_bits_taskID),
    .io_Out_ready(const1_io_Out_ready),
    .io_Out_valid(const1_io_Out_valid),
    .io_Out_bits_taskID(const1_io_Out_bits_taskID)
  );
  ConstFastNode const2 ( // @[bbgemm.scala 253:22]
    .clock(const2_clock),
    .reset(const2_reset),
    .io_enable_ready(const2_io_enable_ready),
    .io_enable_valid(const2_io_enable_valid),
    .io_enable_bits_taskID(const2_io_enable_bits_taskID),
    .io_Out_ready(const2_io_Out_ready),
    .io_Out_valid(const2_io_Out_valid),
    .io_Out_bits_taskID(const2_io_Out_bits_taskID)
  );
  ConstFastNode_3 const3 ( // @[bbgemm.scala 256:22]
    .clock(const3_clock),
    .reset(const3_reset),
    .io_enable_ready(const3_io_enable_ready),
    .io_enable_valid(const3_io_enable_valid),
    .io_Out_ready(const3_io_Out_ready),
    .io_Out_valid(const3_io_Out_valid)
  );
  ConstFastNode const4 ( // @[bbgemm.scala 259:22]
    .clock(const4_clock),
    .reset(const4_reset),
    .io_enable_ready(const4_io_enable_ready),
    .io_enable_valid(const4_io_enable_valid),
    .io_enable_bits_taskID(const4_io_enable_bits_taskID),
    .io_Out_ready(const4_io_Out_ready),
    .io_Out_valid(const4_io_Out_valid),
    .io_Out_bits_taskID(const4_io_Out_bits_taskID)
  );
  ConstFastNode_3 const5 ( // @[bbgemm.scala 262:22]
    .clock(const5_clock),
    .reset(const5_reset),
    .io_enable_ready(const5_io_enable_ready),
    .io_enable_valid(const5_io_enable_valid),
    .io_Out_ready(const5_io_Out_ready),
    .io_Out_valid(const5_io_Out_valid)
  );
  ConstFastNode const6 ( // @[bbgemm.scala 265:22]
    .clock(const6_clock),
    .reset(const6_reset),
    .io_enable_ready(const6_io_enable_ready),
    .io_enable_valid(const6_io_enable_valid),
    .io_enable_bits_taskID(const6_io_enable_bits_taskID),
    .io_Out_ready(const6_io_Out_ready),
    .io_Out_valid(const6_io_Out_valid),
    .io_Out_bits_taskID(const6_io_Out_bits_taskID)
  );
  ConstFastNode_7 const7 ( // @[bbgemm.scala 268:22]
    .clock(const7_clock),
    .reset(const7_reset),
    .io_enable_ready(const7_io_enable_ready),
    .io_enable_valid(const7_io_enable_valid),
    .io_enable_bits_taskID(const7_io_enable_bits_taskID),
    .io_Out_ready(const7_io_Out_ready),
    .io_Out_valid(const7_io_Out_valid),
    .io_Out_bits_taskID(const7_io_Out_bits_taskID)
  );
  ConstFastNode_8 const8 ( // @[bbgemm.scala 271:22]
    .clock(const8_clock),
    .reset(const8_reset),
    .io_enable_ready(const8_io_enable_ready),
    .io_enable_valid(const8_io_enable_valid),
    .io_enable_bits_taskID(const8_io_enable_bits_taskID),
    .io_Out_ready(const8_io_Out_ready),
    .io_Out_valid(const8_io_Out_valid),
    .io_Out_bits_taskID(const8_io_Out_bits_taskID)
  );
  ConstFastNode_7 const9 ( // @[bbgemm.scala 274:22]
    .clock(const9_clock),
    .reset(const9_reset),
    .io_enable_ready(const9_io_enable_ready),
    .io_enable_valid(const9_io_enable_valid),
    .io_enable_bits_taskID(const9_io_enable_bits_taskID),
    .io_Out_ready(const9_io_Out_ready),
    .io_Out_valid(const9_io_Out_valid),
    .io_Out_bits_taskID(const9_io_Out_bits_taskID)
  );
  ConstFastNode_8 const10 ( // @[bbgemm.scala 277:23]
    .clock(const10_clock),
    .reset(const10_reset),
    .io_enable_ready(const10_io_enable_ready),
    .io_enable_valid(const10_io_enable_valid),
    .io_enable_bits_taskID(const10_io_enable_bits_taskID),
    .io_Out_ready(const10_io_Out_ready),
    .io_Out_valid(const10_io_Out_valid),
    .io_Out_bits_taskID(const10_io_Out_bits_taskID)
  );
  ConstFastNode_7 const11 ( // @[bbgemm.scala 280:23]
    .clock(const11_clock),
    .reset(const11_reset),
    .io_enable_ready(const11_io_enable_ready),
    .io_enable_valid(const11_io_enable_valid),
    .io_enable_bits_taskID(const11_io_enable_bits_taskID),
    .io_Out_ready(const11_io_Out_ready),
    .io_Out_valid(const11_io_Out_valid),
    .io_Out_bits_taskID(const11_io_Out_bits_taskID)
  );
  ConstFastNode_12 const12 ( // @[bbgemm.scala 283:23]
    .clock(const12_clock),
    .reset(const12_reset),
    .io_enable_ready(const12_io_enable_ready),
    .io_enable_valid(const12_io_enable_valid),
    .io_enable_bits_taskID(const12_io_enable_bits_taskID),
    .io_Out_ready(const12_io_Out_ready),
    .io_Out_valid(const12_io_Out_valid),
    .io_Out_bits_taskID(const12_io_Out_bits_taskID)
  );
  ConstFastNode_8 const13 ( // @[bbgemm.scala 286:23]
    .clock(const13_clock),
    .reset(const13_reset),
    .io_enable_ready(const13_io_enable_ready),
    .io_enable_valid(const13_io_enable_valid),
    .io_enable_bits_taskID(const13_io_enable_bits_taskID),
    .io_Out_ready(const13_io_Out_ready),
    .io_Out_valid(const13_io_Out_valid),
    .io_Out_bits_taskID(const13_io_Out_bits_taskID)
  );
  ConstFastNode_12 const14 ( // @[bbgemm.scala 289:23]
    .clock(const14_clock),
    .reset(const14_reset),
    .io_enable_ready(const14_io_enable_ready),
    .io_enable_valid(const14_io_enable_valid),
    .io_enable_bits_taskID(const14_io_enable_bits_taskID),
    .io_Out_ready(const14_io_Out_ready),
    .io_Out_valid(const14_io_Out_valid),
    .io_Out_bits_taskID(const14_io_Out_bits_taskID)
  );
  ConstFastNode_8 const15 ( // @[bbgemm.scala 292:23]
    .clock(const15_clock),
    .reset(const15_reset),
    .io_enable_ready(const15_io_enable_ready),
    .io_enable_valid(const15_io_enable_valid),
    .io_enable_bits_taskID(const15_io_enable_bits_taskID),
    .io_Out_ready(const15_io_Out_ready),
    .io_Out_valid(const15_io_Out_valid),
    .io_Out_bits_taskID(const15_io_Out_bits_taskID)
  );
  ConstFastNode_12 const16 ( // @[bbgemm.scala 295:23]
    .clock(const16_clock),
    .reset(const16_reset),
    .io_enable_ready(const16_io_enable_ready),
    .io_enable_valid(const16_io_enable_valid),
    .io_enable_bits_taskID(const16_io_enable_bits_taskID),
    .io_Out_ready(const16_io_Out_ready),
    .io_Out_valid(const16_io_Out_valid),
    .io_Out_bits_taskID(const16_io_Out_bits_taskID)
  );
  assign io_in_ready = InputSplitter_io_In_ready; // @[bbgemm.scala 54:23]
  assign io_MemReq_valid = MemCtrl_io_MemReq_valid; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_addr = MemCtrl_io_MemReq_bits_addr; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_data = MemCtrl_io_MemReq_bits_data; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_mask = MemCtrl_io_MemReq_bits_mask; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_tag = MemCtrl_io_MemReq_bits_tag; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_taskID = MemCtrl_io_MemReq_bits_taskID; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_iswrite = MemCtrl_io_MemReq_bits_iswrite; // @[bbgemm.scala 50:13]
  assign io_MemReq_bits_tile = 32'h0; // @[bbgemm.scala 50:13]
  assign io_out_valid = ret_43_io_Out_valid; // @[bbgemm.scala 855:10]
  assign io_out_bits_enable_taskID = ret_43_io_Out_bits_enable_taskID; // @[bbgemm.scala 855:10]
  assign io_out_bits_enable_control = ret_43_io_Out_bits_enable_control; // @[bbgemm.scala 855:10]
  assign MemCtrl_clock = clock;
  assign MemCtrl_reset = reset;
  assign MemCtrl_io_WriteIn_0_valid = st_27_io_memReq_valid; // @[bbgemm.scala 727:25]
  assign MemCtrl_io_WriteIn_0_bits_address = st_27_io_memReq_bits_address; // @[bbgemm.scala 727:25]
  assign MemCtrl_io_WriteIn_0_bits_data = st_27_io_memReq_bits_data; // @[bbgemm.scala 727:25]
  assign MemCtrl_io_WriteIn_0_bits_taskID = st_27_io_memReq_bits_taskID; // @[bbgemm.scala 727:25]
  assign MemCtrl_io_ReadIn_0_valid = ld_14_io_memReq_valid; // @[bbgemm.scala 715:24]
  assign MemCtrl_io_ReadIn_0_bits_address = ld_14_io_memReq_bits_address; // @[bbgemm.scala 715:24]
  assign MemCtrl_io_ReadIn_0_bits_taskID = ld_14_io_memReq_bits_taskID; // @[bbgemm.scala 715:24]
  assign MemCtrl_io_ReadIn_1_valid = ld_20_io_memReq_valid; // @[bbgemm.scala 719:24]
  assign MemCtrl_io_ReadIn_1_bits_address = ld_20_io_memReq_bits_address; // @[bbgemm.scala 719:24]
  assign MemCtrl_io_ReadIn_1_bits_taskID = ld_20_io_memReq_bits_taskID; // @[bbgemm.scala 719:24]
  assign MemCtrl_io_ReadIn_2_valid = ld_25_io_memReq_valid; // @[bbgemm.scala 723:24]
  assign MemCtrl_io_ReadIn_2_bits_address = ld_25_io_memReq_bits_address; // @[bbgemm.scala 723:24]
  assign MemCtrl_io_ReadIn_2_bits_taskID = ld_25_io_memReq_bits_taskID; // @[bbgemm.scala 723:24]
  assign MemCtrl_io_MemResp_valid = io_MemResp_valid; // @[bbgemm.scala 51:22]
  assign MemCtrl_io_MemResp_bits_data = io_MemResp_bits_data; // @[bbgemm.scala 51:22]
  assign MemCtrl_io_MemResp_bits_tag = io_MemResp_bits_tag; // @[bbgemm.scala 51:22]
  assign MemCtrl_io_MemResp_bits_iswrite = io_MemResp_bits_iswrite; // @[bbgemm.scala 51:22]
  assign MemCtrl_io_MemReq_ready = io_MemReq_ready; // @[bbgemm.scala 50:13]
  assign InputSplitter_clock = clock;
  assign InputSplitter_reset = reset;
  assign InputSplitter_io_In_valid = io_in_valid; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_enable_taskID = io_in_bits_enable_taskID; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_enable_control = io_in_bits_enable_control; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_data_field2_taskID = io_in_bits_data_field2_taskID; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_data_field2_data = io_in_bits_data_field2_data; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_taskID = io_in_bits_data_field1_taskID; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_data = io_in_bits_data_field1_data; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_data_field0_taskID = io_in_bits_data_field0_taskID; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_In_bits_data_field0_data = io_in_bits_data_field0_data; // @[bbgemm.scala 54:23]
  assign InputSplitter_io_Out_enable_ready = bb_0_io_predicateIn_0_ready; // @[bbgemm.scala 303:26]
  assign InputSplitter_io_Out_data_field2_0_ready = Loop_4_io_InLiveIn_2_ready; // @[bbgemm.scala 441:25]
  assign InputSplitter_io_Out_data_field1_0_ready = Loop_4_io_InLiveIn_1_ready; // @[bbgemm.scala 439:25]
  assign InputSplitter_io_Out_data_field0_0_ready = Loop_4_io_InLiveIn_0_ready; // @[bbgemm.scala 437:25]
  assign Loop_0_clock = clock;
  assign Loop_0_reset = reset;
  assign Loop_0_io_enable_valid = br_15_io_Out_0_valid; // @[bbgemm.scala 353:20]
  assign Loop_0_io_enable_bits_taskID = br_15_io_Out_0_bits_taskID; // @[bbgemm.scala 353:20]
  assign Loop_0_io_enable_bits_control = br_15_io_Out_0_bits_control; // @[bbgemm.scala 353:20]
  assign Loop_0_io_InLiveIn_0_valid = binaryOp_10_io_Out_0_valid; // @[bbgemm.scala 395:25]
  assign Loop_0_io_InLiveIn_0_bits_data = binaryOp_10_io_Out_0_bits_data; // @[bbgemm.scala 395:25]
  assign Loop_0_io_InLiveIn_1_valid = ld_14_io_Out_0_valid; // @[bbgemm.scala 397:25]
  assign Loop_0_io_InLiveIn_1_bits_taskID = ld_14_io_Out_0_bits_taskID; // @[bbgemm.scala 397:25]
  assign Loop_0_io_InLiveIn_1_bits_data = ld_14_io_Out_0_bits_data; // @[bbgemm.scala 397:25]
  assign Loop_0_io_InLiveIn_2_valid = Loop_1_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 399:25]
  assign Loop_0_io_InLiveIn_2_bits_data = Loop_1_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 399:25]
  assign Loop_0_io_InLiveIn_3_valid = Loop_1_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 401:25]
  assign Loop_0_io_InLiveIn_3_bits_taskID = Loop_1_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 401:25]
  assign Loop_0_io_InLiveIn_3_bits_data = Loop_1_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 401:25]
  assign Loop_0_io_InLiveIn_4_valid = Loop_1_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 403:25]
  assign Loop_0_io_InLiveIn_4_bits_taskID = Loop_1_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 403:25]
  assign Loop_0_io_InLiveIn_4_bits_data = Loop_1_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 403:25]
  assign Loop_0_io_InLiveIn_5_valid = Loop_1_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 405:25]
  assign Loop_0_io_InLiveIn_5_bits_data = Loop_1_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 405:25]
  assign Loop_0_io_OutLiveIn_field5_0_ready = binaryOp_17_io_RightIO_ready; // @[bbgemm.scala 459:26]
  assign Loop_0_io_OutLiveIn_field5_1_ready = binaryOp_22_io_RightIO_ready; // @[bbgemm.scala 461:26]
  assign Loop_0_io_OutLiveIn_field4_0_ready = Gep_19_io_baseAddress_ready; // @[bbgemm.scala 457:25]
  assign Loop_0_io_OutLiveIn_field3_0_ready = Gep_24_io_baseAddress_ready; // @[bbgemm.scala 455:25]
  assign Loop_0_io_OutLiveIn_field2_0_ready = binaryOp_23_io_RightIO_ready; // @[bbgemm.scala 453:26]
  assign Loop_0_io_OutLiveIn_field1_0_ready = FP_21_io_LeftIO_ready; // @[bbgemm.scala 451:19]
  assign Loop_0_io_OutLiveIn_field0_0_ready = binaryOp_18_io_RightIO_ready; // @[bbgemm.scala 449:26]
  assign Loop_0_io_activate_loop_start_ready = bb_5_io_predicateIn_1_ready; // @[bbgemm.scala 327:26]
  assign Loop_0_io_activate_loop_back_ready = bb_5_io_predicateIn_0_ready; // @[bbgemm.scala 329:26]
  assign Loop_0_io_loopBack_0_valid = br_30_io_FalseOutput_0_valid; // @[bbgemm.scala 355:25]
  assign Loop_0_io_loopBack_0_bits_taskID = br_30_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 355:25]
  assign Loop_0_io_loopBack_0_bits_control = br_30_io_FalseOutput_0_bits_control; // @[bbgemm.scala 355:25]
  assign Loop_0_io_loopFinish_0_valid = br_30_io_TrueOutput_0_valid; // @[bbgemm.scala 357:27]
  assign Loop_0_io_loopFinish_0_bits_control = br_30_io_TrueOutput_0_bits_control; // @[bbgemm.scala 357:27]
  assign Loop_0_io_CarryDepenIn_0_valid = binaryOp_28_io_Out_0_valid; // @[bbgemm.scala 489:29]
  assign Loop_0_io_CarryDepenIn_0_bits_taskID = binaryOp_28_io_Out_0_bits_taskID; // @[bbgemm.scala 489:29]
  assign Loop_0_io_CarryDepenIn_0_bits_data = binaryOp_28_io_Out_0_bits_data; // @[bbgemm.scala 489:29]
  assign Loop_0_io_CarryDepenOut_field0_0_ready = phi16_io_InData_1_ready; // @[bbgemm.scala 505:22]
  assign Loop_0_io_loopExit_0_ready = bb_6_io_predicateIn_0_ready; // @[bbgemm.scala 331:26]
  assign Loop_1_clock = clock;
  assign Loop_1_reset = reset;
  assign Loop_1_io_enable_valid = br_7_io_Out_0_valid; // @[bbgemm.scala 359:20]
  assign Loop_1_io_enable_bits_taskID = br_7_io_Out_0_bits_taskID; // @[bbgemm.scala 359:20]
  assign Loop_1_io_enable_bits_control = br_7_io_Out_0_bits_control; // @[bbgemm.scala 359:20]
  assign Loop_1_io_InLiveIn_0_valid = binaryOp_6_io_Out_0_valid; // @[bbgemm.scala 407:25]
  assign Loop_1_io_InLiveIn_0_bits_data = binaryOp_6_io_Out_0_bits_data; // @[bbgemm.scala 407:25]
  assign Loop_1_io_InLiveIn_1_valid = Loop_2_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 409:25]
  assign Loop_1_io_InLiveIn_1_bits_taskID = Loop_2_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 409:25]
  assign Loop_1_io_InLiveIn_1_bits_data = Loop_2_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 409:25]
  assign Loop_1_io_InLiveIn_2_valid = Loop_2_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 411:25]
  assign Loop_1_io_InLiveIn_2_bits_taskID = Loop_2_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 411:25]
  assign Loop_1_io_InLiveIn_2_bits_data = Loop_2_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 411:25]
  assign Loop_1_io_InLiveIn_3_valid = Loop_2_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 413:25]
  assign Loop_1_io_InLiveIn_3_bits_data = Loop_2_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 413:25]
  assign Loop_1_io_InLiveIn_4_valid = Loop_2_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 415:25]
  assign Loop_1_io_InLiveIn_4_bits_data = Loop_2_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 415:25]
  assign Loop_1_io_InLiveIn_5_valid = Loop_2_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 417:25]
  assign Loop_1_io_InLiveIn_5_bits_taskID = Loop_2_io_OutLiveIn_field3_0_bits_taskID; // @[bbgemm.scala 417:25]
  assign Loop_1_io_InLiveIn_5_bits_data = Loop_2_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 417:25]
  assign Loop_1_io_OutLiveIn_field5_0_ready = Gep_13_io_baseAddress_ready; // @[bbgemm.scala 469:25]
  assign Loop_1_io_OutLiveIn_field4_0_ready = binaryOp_9_io_RightIO_ready; // @[bbgemm.scala 465:25]
  assign Loop_1_io_OutLiveIn_field4_1_ready = binaryOp_11_io_RightIO_ready; // @[bbgemm.scala 467:26]
  assign Loop_1_io_OutLiveIn_field3_0_ready = Loop_0_io_InLiveIn_5_ready; // @[bbgemm.scala 405:25]
  assign Loop_1_io_OutLiveIn_field2_0_ready = Loop_0_io_InLiveIn_4_ready; // @[bbgemm.scala 403:25]
  assign Loop_1_io_OutLiveIn_field1_0_ready = Loop_0_io_InLiveIn_3_ready; // @[bbgemm.scala 401:25]
  assign Loop_1_io_OutLiveIn_field0_0_ready = Loop_0_io_InLiveIn_2_ready; // @[bbgemm.scala 399:25]
  assign Loop_1_io_OutLiveIn_field0_1_ready = binaryOp_12_io_RightIO_ready; // @[bbgemm.scala 463:26]
  assign Loop_1_io_activate_loop_start_ready = bb_4_io_predicateIn_1_ready; // @[bbgemm.scala 323:26]
  assign Loop_1_io_activate_loop_back_ready = bb_4_io_predicateIn_0_ready; // @[bbgemm.scala 325:26]
  assign Loop_1_io_loopBack_0_valid = br_33_io_FalseOutput_0_valid; // @[bbgemm.scala 361:25]
  assign Loop_1_io_loopBack_0_bits_taskID = br_33_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 361:25]
  assign Loop_1_io_loopBack_0_bits_control = br_33_io_FalseOutput_0_bits_control; // @[bbgemm.scala 361:25]
  assign Loop_1_io_loopFinish_0_valid = br_33_io_TrueOutput_0_valid; // @[bbgemm.scala 363:27]
  assign Loop_1_io_loopFinish_0_bits_control = br_33_io_TrueOutput_0_bits_control; // @[bbgemm.scala 363:27]
  assign Loop_1_io_CarryDepenIn_0_valid = binaryOp_31_io_Out_0_valid; // @[bbgemm.scala 491:29]
  assign Loop_1_io_CarryDepenIn_0_bits_taskID = binaryOp_31_io_Out_0_bits_taskID; // @[bbgemm.scala 491:29]
  assign Loop_1_io_CarryDepenIn_0_bits_data = binaryOp_31_io_Out_0_bits_data; // @[bbgemm.scala 491:29]
  assign Loop_1_io_CarryDepenOut_field0_0_ready = phi8_io_InData_1_ready; // @[bbgemm.scala 507:21]
  assign Loop_1_io_loopExit_0_ready = bb_7_io_predicateIn_0_ready; // @[bbgemm.scala 333:26]
  assign Loop_2_clock = clock;
  assign Loop_2_reset = reset;
  assign Loop_2_io_enable_valid = br_4_io_Out_0_valid; // @[bbgemm.scala 365:20]
  assign Loop_2_io_enable_bits_taskID = br_4_io_Out_0_bits_taskID; // @[bbgemm.scala 365:20]
  assign Loop_2_io_enable_bits_control = br_4_io_Out_0_bits_control; // @[bbgemm.scala 365:20]
  assign Loop_2_io_InLiveIn_0_valid = phi3_io_Out_0_valid; // @[bbgemm.scala 419:25]
  assign Loop_2_io_InLiveIn_0_bits_data = phi3_io_Out_0_bits_data; // @[bbgemm.scala 419:25]
  assign Loop_2_io_InLiveIn_1_valid = Loop_3_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 421:25]
  assign Loop_2_io_InLiveIn_1_bits_taskID = Loop_3_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 421:25]
  assign Loop_2_io_InLiveIn_1_bits_data = Loop_3_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 421:25]
  assign Loop_2_io_InLiveIn_2_valid = Loop_3_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 423:25]
  assign Loop_2_io_InLiveIn_2_bits_taskID = Loop_3_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 423:25]
  assign Loop_2_io_InLiveIn_2_bits_data = Loop_3_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 423:25]
  assign Loop_2_io_InLiveIn_3_valid = Loop_3_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 425:25]
  assign Loop_2_io_InLiveIn_3_bits_taskID = Loop_3_io_OutLiveIn_field3_0_bits_taskID; // @[bbgemm.scala 425:25]
  assign Loop_2_io_InLiveIn_3_bits_data = Loop_3_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 425:25]
  assign Loop_2_io_InLiveIn_4_valid = Loop_3_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 427:25]
  assign Loop_2_io_InLiveIn_4_bits_data = Loop_3_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 427:25]
  assign Loop_2_io_OutLiveIn_field4_0_ready = Loop_1_io_InLiveIn_3_ready; // @[bbgemm.scala 413:25]
  assign Loop_2_io_OutLiveIn_field3_0_ready = Loop_1_io_InLiveIn_5_ready; // @[bbgemm.scala 417:25]
  assign Loop_2_io_OutLiveIn_field2_0_ready = Loop_1_io_InLiveIn_2_ready; // @[bbgemm.scala 411:25]
  assign Loop_2_io_OutLiveIn_field1_0_ready = Loop_1_io_InLiveIn_1_ready; // @[bbgemm.scala 409:25]
  assign Loop_2_io_OutLiveIn_field0_0_ready = Loop_1_io_InLiveIn_4_ready; // @[bbgemm.scala 415:25]
  assign Loop_2_io_activate_loop_start_ready = bb_3_io_predicateIn_1_ready; // @[bbgemm.scala 319:26]
  assign Loop_2_io_activate_loop_back_ready = bb_3_io_predicateIn_0_ready; // @[bbgemm.scala 321:26]
  assign Loop_2_io_loopBack_0_valid = br_36_io_FalseOutput_0_valid; // @[bbgemm.scala 367:25]
  assign Loop_2_io_loopBack_0_bits_taskID = br_36_io_FalseOutput_0_bits_taskID; // @[bbgemm.scala 367:25]
  assign Loop_2_io_loopBack_0_bits_control = br_36_io_FalseOutput_0_bits_control; // @[bbgemm.scala 367:25]
  assign Loop_2_io_loopFinish_0_valid = br_36_io_TrueOutput_0_valid; // @[bbgemm.scala 369:27]
  assign Loop_2_io_loopFinish_0_bits_control = br_36_io_TrueOutput_0_bits_control; // @[bbgemm.scala 369:27]
  assign Loop_2_io_CarryDepenIn_0_valid = binaryOp_34_io_Out_0_valid; // @[bbgemm.scala 493:29]
  assign Loop_2_io_CarryDepenIn_0_bits_taskID = binaryOp_34_io_Out_0_bits_taskID; // @[bbgemm.scala 493:29]
  assign Loop_2_io_CarryDepenIn_0_bits_data = binaryOp_34_io_Out_0_bits_data; // @[bbgemm.scala 493:29]
  assign Loop_2_io_CarryDepenOut_field0_0_ready = phi5_io_InData_1_ready; // @[bbgemm.scala 509:21]
  assign Loop_2_io_loopExit_0_ready = bb_8_io_predicateIn_0_ready; // @[bbgemm.scala 335:26]
  assign Loop_3_clock = clock;
  assign Loop_3_reset = reset;
  assign Loop_3_io_enable_valid = br_2_io_Out_0_valid; // @[bbgemm.scala 371:20]
  assign Loop_3_io_enable_bits_taskID = br_2_io_Out_0_bits_taskID; // @[bbgemm.scala 371:20]
  assign Loop_3_io_enable_bits_control = br_2_io_Out_0_bits_control; // @[bbgemm.scala 371:20]
  assign Loop_3_io_InLiveIn_0_valid = phi1_io_Out_0_valid; // @[bbgemm.scala 429:25]
  assign Loop_3_io_InLiveIn_0_bits_data = phi1_io_Out_0_bits_data; // @[bbgemm.scala 429:25]
  assign Loop_3_io_InLiveIn_1_valid = Loop_4_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 431:25]
  assign Loop_3_io_InLiveIn_1_bits_taskID = Loop_4_io_OutLiveIn_field2_0_bits_taskID; // @[bbgemm.scala 431:25]
  assign Loop_3_io_InLiveIn_1_bits_data = Loop_4_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 431:25]
  assign Loop_3_io_InLiveIn_2_valid = Loop_4_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 433:25]
  assign Loop_3_io_InLiveIn_2_bits_taskID = Loop_4_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 433:25]
  assign Loop_3_io_InLiveIn_2_bits_data = Loop_4_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 433:25]
  assign Loop_3_io_InLiveIn_3_valid = Loop_4_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 435:25]
  assign Loop_3_io_InLiveIn_3_bits_taskID = Loop_4_io_OutLiveIn_field0_0_bits_taskID; // @[bbgemm.scala 435:25]
  assign Loop_3_io_InLiveIn_3_bits_data = Loop_4_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 435:25]
  assign Loop_3_io_OutLiveIn_field3_0_ready = Loop_2_io_InLiveIn_3_ready; // @[bbgemm.scala 425:25]
  assign Loop_3_io_OutLiveIn_field2_0_ready = Loop_2_io_InLiveIn_2_ready; // @[bbgemm.scala 423:25]
  assign Loop_3_io_OutLiveIn_field1_0_ready = Loop_2_io_InLiveIn_1_ready; // @[bbgemm.scala 421:25]
  assign Loop_3_io_OutLiveIn_field0_0_ready = Loop_2_io_InLiveIn_4_ready; // @[bbgemm.scala 427:25]
  assign Loop_3_io_activate_loop_start_ready = bb_2_io_predicateIn_0_ready; // @[bbgemm.scala 315:26]
  assign Loop_3_io_activate_loop_back_ready = bb_2_io_predicateIn_1_ready; // @[bbgemm.scala 317:26]
  assign Loop_3_io_loopBack_0_valid = br_39_io_TrueOutput_0_valid; // @[bbgemm.scala 373:25]
  assign Loop_3_io_loopBack_0_bits_taskID = br_39_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 373:25]
  assign Loop_3_io_loopBack_0_bits_control = br_39_io_TrueOutput_0_bits_control; // @[bbgemm.scala 373:25]
  assign Loop_3_io_loopFinish_0_valid = br_39_io_FalseOutput_0_valid; // @[bbgemm.scala 375:27]
  assign Loop_3_io_loopFinish_0_bits_control = br_39_io_FalseOutput_0_bits_control; // @[bbgemm.scala 375:27]
  assign Loop_3_io_CarryDepenIn_0_valid = binaryOp_37_io_Out_0_valid; // @[bbgemm.scala 495:29]
  assign Loop_3_io_CarryDepenIn_0_bits_taskID = binaryOp_37_io_Out_0_bits_taskID; // @[bbgemm.scala 495:29]
  assign Loop_3_io_CarryDepenIn_0_bits_data = binaryOp_37_io_Out_0_bits_data; // @[bbgemm.scala 495:29]
  assign Loop_3_io_CarryDepenOut_field0_0_ready = phi3_io_InData_1_ready; // @[bbgemm.scala 511:21]
  assign Loop_3_io_loopExit_0_ready = bb_9_io_predicateIn_0_ready; // @[bbgemm.scala 337:26]
  assign Loop_4_clock = clock;
  assign Loop_4_reset = reset;
  assign Loop_4_io_enable_valid = br_0_io_Out_0_valid; // @[bbgemm.scala 377:20]
  assign Loop_4_io_enable_bits_taskID = br_0_io_Out_0_bits_taskID; // @[bbgemm.scala 377:20]
  assign Loop_4_io_enable_bits_control = br_0_io_Out_0_bits_control; // @[bbgemm.scala 377:20]
  assign Loop_4_io_InLiveIn_0_valid = InputSplitter_io_Out_data_field0_0_valid; // @[bbgemm.scala 437:25]
  assign Loop_4_io_InLiveIn_0_bits_taskID = InputSplitter_io_Out_data_field0_0_bits_taskID; // @[bbgemm.scala 437:25]
  assign Loop_4_io_InLiveIn_0_bits_data = InputSplitter_io_Out_data_field0_0_bits_data; // @[bbgemm.scala 437:25]
  assign Loop_4_io_InLiveIn_1_valid = InputSplitter_io_Out_data_field1_0_valid; // @[bbgemm.scala 439:25]
  assign Loop_4_io_InLiveIn_1_bits_taskID = InputSplitter_io_Out_data_field1_0_bits_taskID; // @[bbgemm.scala 439:25]
  assign Loop_4_io_InLiveIn_1_bits_data = InputSplitter_io_Out_data_field1_0_bits_data; // @[bbgemm.scala 439:25]
  assign Loop_4_io_InLiveIn_2_valid = InputSplitter_io_Out_data_field2_0_valid; // @[bbgemm.scala 441:25]
  assign Loop_4_io_InLiveIn_2_bits_taskID = InputSplitter_io_Out_data_field2_0_bits_taskID; // @[bbgemm.scala 441:25]
  assign Loop_4_io_InLiveIn_2_bits_data = InputSplitter_io_Out_data_field2_0_bits_data; // @[bbgemm.scala 441:25]
  assign Loop_4_io_OutLiveIn_field2_0_ready = Loop_3_io_InLiveIn_1_ready; // @[bbgemm.scala 431:25]
  assign Loop_4_io_OutLiveIn_field1_0_ready = Loop_3_io_InLiveIn_2_ready; // @[bbgemm.scala 433:25]
  assign Loop_4_io_OutLiveIn_field0_0_ready = Loop_3_io_InLiveIn_3_ready; // @[bbgemm.scala 435:25]
  assign Loop_4_io_activate_loop_start_ready = bb_1_io_predicateIn_0_ready; // @[bbgemm.scala 311:26]
  assign Loop_4_io_activate_loop_back_ready = bb_1_io_predicateIn_1_ready; // @[bbgemm.scala 313:26]
  assign Loop_4_io_loopBack_0_valid = br_42_io_TrueOutput_0_valid; // @[bbgemm.scala 379:25]
  assign Loop_4_io_loopBack_0_bits_taskID = br_42_io_TrueOutput_0_bits_taskID; // @[bbgemm.scala 379:25]
  assign Loop_4_io_loopBack_0_bits_control = br_42_io_TrueOutput_0_bits_control; // @[bbgemm.scala 379:25]
  assign Loop_4_io_loopFinish_0_valid = br_42_io_FalseOutput_0_valid; // @[bbgemm.scala 381:27]
  assign Loop_4_io_loopFinish_0_bits_control = br_42_io_FalseOutput_0_bits_control; // @[bbgemm.scala 381:27]
  assign Loop_4_io_CarryDepenIn_0_valid = binaryOp_40_io_Out_0_valid; // @[bbgemm.scala 497:29]
  assign Loop_4_io_CarryDepenIn_0_bits_taskID = binaryOp_40_io_Out_0_bits_taskID; // @[bbgemm.scala 497:29]
  assign Loop_4_io_CarryDepenIn_0_bits_data = binaryOp_40_io_Out_0_bits_data; // @[bbgemm.scala 497:29]
  assign Loop_4_io_CarryDepenOut_field0_0_ready = phi1_io_InData_1_ready; // @[bbgemm.scala 513:21]
  assign Loop_4_io_loopExit_0_ready = bb_10_io_predicateIn_0_ready; // @[bbgemm.scala 339:27]
  assign bb_0_clock = clock;
  assign bb_0_reset = reset;
  assign bb_0_io_predicateIn_0_valid = InputSplitter_io_Out_enable_valid; // @[bbgemm.scala 303:26]
  assign bb_0_io_predicateIn_0_bits_taskID = InputSplitter_io_Out_enable_bits_taskID; // @[bbgemm.scala 303:26]
  assign bb_0_io_predicateIn_0_bits_control = InputSplitter_io_Out_enable_bits_control; // @[bbgemm.scala 303:26]
  assign bb_0_io_Out_0_ready = br_0_io_enable_ready; // @[bbgemm.scala 521:18]
  assign bb_1_clock = clock;
  assign bb_1_reset = reset;
  assign bb_1_io_MaskBB_0_ready = phi1_io_Mask_ready; // @[bbgemm.scala 693:16]
  assign bb_1_io_Out_0_ready = const0_io_enable_ready; // @[bbgemm.scala 524:20]
  assign bb_1_io_Out_1_ready = phi1_io_enable_ready; // @[bbgemm.scala 526:18]
  assign bb_1_io_Out_2_ready = br_2_io_enable_ready; // @[bbgemm.scala 529:18]
  assign bb_1_io_predicateIn_0_valid = Loop_4_io_activate_loop_start_valid; // @[bbgemm.scala 311:26]
  assign bb_1_io_predicateIn_0_bits_taskID = Loop_4_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 311:26]
  assign bb_1_io_predicateIn_0_bits_control = Loop_4_io_activate_loop_start_bits_control; // @[bbgemm.scala 311:26]
  assign bb_1_io_predicateIn_1_valid = Loop_4_io_activate_loop_back_valid; // @[bbgemm.scala 313:26]
  assign bb_1_io_predicateIn_1_bits_taskID = Loop_4_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 313:26]
  assign bb_1_io_predicateIn_1_bits_control = Loop_4_io_activate_loop_back_bits_control; // @[bbgemm.scala 313:26]
  assign bb_2_clock = clock;
  assign bb_2_reset = reset;
  assign bb_2_io_MaskBB_0_ready = phi3_io_Mask_ready; // @[bbgemm.scala 695:16]
  assign bb_2_io_Out_0_ready = const1_io_enable_ready; // @[bbgemm.scala 532:20]
  assign bb_2_io_Out_1_ready = phi3_io_enable_ready; // @[bbgemm.scala 534:18]
  assign bb_2_io_Out_2_ready = br_4_io_enable_ready; // @[bbgemm.scala 537:18]
  assign bb_2_io_predicateIn_0_valid = Loop_3_io_activate_loop_start_valid; // @[bbgemm.scala 315:26]
  assign bb_2_io_predicateIn_0_bits_taskID = Loop_3_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 315:26]
  assign bb_2_io_predicateIn_0_bits_control = Loop_3_io_activate_loop_start_bits_control; // @[bbgemm.scala 315:26]
  assign bb_2_io_predicateIn_1_valid = Loop_3_io_activate_loop_back_valid; // @[bbgemm.scala 317:26]
  assign bb_2_io_predicateIn_1_bits_taskID = Loop_3_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 317:26]
  assign bb_2_io_predicateIn_1_bits_control = Loop_3_io_activate_loop_back_bits_control; // @[bbgemm.scala 317:26]
  assign bb_3_clock = clock;
  assign bb_3_reset = reset;
  assign bb_3_io_MaskBB_0_ready = phi5_io_Mask_ready; // @[bbgemm.scala 697:16]
  assign bb_3_io_Out_0_ready = const2_io_enable_ready; // @[bbgemm.scala 540:20]
  assign bb_3_io_Out_1_ready = const3_io_enable_ready; // @[bbgemm.scala 542:20]
  assign bb_3_io_Out_2_ready = phi5_io_enable_ready; // @[bbgemm.scala 544:18]
  assign bb_3_io_Out_3_ready = binaryOp_6_io_enable_ready; // @[bbgemm.scala 547:24]
  assign bb_3_io_Out_4_ready = br_7_io_enable_ready; // @[bbgemm.scala 550:18]
  assign bb_3_io_predicateIn_0_valid = Loop_2_io_activate_loop_back_valid; // @[bbgemm.scala 321:26]
  assign bb_3_io_predicateIn_0_bits_taskID = Loop_2_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 321:26]
  assign bb_3_io_predicateIn_0_bits_control = Loop_2_io_activate_loop_back_bits_control; // @[bbgemm.scala 321:26]
  assign bb_3_io_predicateIn_1_valid = Loop_2_io_activate_loop_start_valid; // @[bbgemm.scala 319:26]
  assign bb_3_io_predicateIn_1_bits_taskID = Loop_2_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 319:26]
  assign bb_3_io_predicateIn_1_bits_control = Loop_2_io_activate_loop_start_bits_control; // @[bbgemm.scala 319:26]
  assign bb_4_clock = clock;
  assign bb_4_reset = reset;
  assign bb_4_io_MaskBB_0_ready = phi8_io_Mask_ready; // @[bbgemm.scala 699:16]
  assign bb_4_io_Out_0_ready = const4_io_enable_ready; // @[bbgemm.scala 553:20]
  assign bb_4_io_Out_1_ready = const5_io_enable_ready; // @[bbgemm.scala 555:20]
  assign bb_4_io_Out_2_ready = phi8_io_enable_ready; // @[bbgemm.scala 557:18]
  assign bb_4_io_Out_3_ready = binaryOp_9_io_enable_ready; // @[bbgemm.scala 560:24]
  assign bb_4_io_Out_4_ready = binaryOp_10_io_enable_ready; // @[bbgemm.scala 563:25]
  assign bb_4_io_Out_5_ready = binaryOp_11_io_enable_ready; // @[bbgemm.scala 566:25]
  assign bb_4_io_Out_6_ready = binaryOp_12_io_enable_ready; // @[bbgemm.scala 569:25]
  assign bb_4_io_Out_7_ready = Gep_13_io_enable_ready; // @[bbgemm.scala 572:20]
  assign bb_4_io_Out_8_ready = ld_14_io_enable_ready; // @[bbgemm.scala 575:19]
  assign bb_4_io_Out_9_ready = br_15_io_enable_ready; // @[bbgemm.scala 578:19]
  assign bb_4_io_predicateIn_0_valid = Loop_1_io_activate_loop_back_valid; // @[bbgemm.scala 325:26]
  assign bb_4_io_predicateIn_0_bits_taskID = Loop_1_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 325:26]
  assign bb_4_io_predicateIn_0_bits_control = Loop_1_io_activate_loop_back_bits_control; // @[bbgemm.scala 325:26]
  assign bb_4_io_predicateIn_1_valid = Loop_1_io_activate_loop_start_valid; // @[bbgemm.scala 323:26]
  assign bb_4_io_predicateIn_1_bits_taskID = Loop_1_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 323:26]
  assign bb_4_io_predicateIn_1_bits_control = Loop_1_io_activate_loop_start_bits_control; // @[bbgemm.scala 323:26]
  assign bb_5_clock = clock;
  assign bb_5_reset = reset;
  assign bb_5_io_MaskBB_0_ready = phi16_io_Mask_ready; // @[bbgemm.scala 701:17]
  assign bb_5_io_Out_0_ready = const6_io_enable_ready; // @[bbgemm.scala 581:20]
  assign bb_5_io_Out_1_ready = const7_io_enable_ready; // @[bbgemm.scala 583:20]
  assign bb_5_io_Out_2_ready = const8_io_enable_ready; // @[bbgemm.scala 585:20]
  assign bb_5_io_Out_3_ready = phi16_io_enable_ready; // @[bbgemm.scala 587:19]
  assign bb_5_io_Out_4_ready = binaryOp_17_io_enable_ready; // @[bbgemm.scala 590:25]
  assign bb_5_io_Out_5_ready = binaryOp_18_io_enable_ready; // @[bbgemm.scala 593:25]
  assign bb_5_io_Out_6_ready = Gep_19_io_enable_ready; // @[bbgemm.scala 596:20]
  assign bb_5_io_Out_7_ready = ld_20_io_enable_ready; // @[bbgemm.scala 599:19]
  assign bb_5_io_Out_8_ready = FP_21_io_enable_ready; // @[bbgemm.scala 602:19]
  assign bb_5_io_Out_9_ready = binaryOp_22_io_enable_ready; // @[bbgemm.scala 605:25]
  assign bb_5_io_Out_10_ready = binaryOp_23_io_enable_ready; // @[bbgemm.scala 608:25]
  assign bb_5_io_Out_11_ready = Gep_24_io_enable_ready; // @[bbgemm.scala 611:20]
  assign bb_5_io_Out_12_ready = ld_25_io_enable_ready; // @[bbgemm.scala 614:19]
  assign bb_5_io_Out_13_ready = FP_26_io_enable_ready; // @[bbgemm.scala 617:19]
  assign bb_5_io_Out_14_ready = st_27_io_enable_ready; // @[bbgemm.scala 620:19]
  assign bb_5_io_Out_15_ready = binaryOp_28_io_enable_ready; // @[bbgemm.scala 623:25]
  assign bb_5_io_Out_16_ready = icmp_29_io_enable_ready; // @[bbgemm.scala 626:21]
  assign bb_5_io_Out_17_ready = br_30_io_enable_ready; // @[bbgemm.scala 629:19]
  assign bb_5_io_predicateIn_0_valid = Loop_0_io_activate_loop_back_valid; // @[bbgemm.scala 329:26]
  assign bb_5_io_predicateIn_0_bits_taskID = Loop_0_io_activate_loop_back_bits_taskID; // @[bbgemm.scala 329:26]
  assign bb_5_io_predicateIn_0_bits_control = Loop_0_io_activate_loop_back_bits_control; // @[bbgemm.scala 329:26]
  assign bb_5_io_predicateIn_1_valid = Loop_0_io_activate_loop_start_valid; // @[bbgemm.scala 327:26]
  assign bb_5_io_predicateIn_1_bits_taskID = Loop_0_io_activate_loop_start_bits_taskID; // @[bbgemm.scala 327:26]
  assign bb_5_io_predicateIn_1_bits_control = Loop_0_io_activate_loop_start_bits_control; // @[bbgemm.scala 327:26]
  assign bb_6_clock = clock;
  assign bb_6_reset = reset;
  assign bb_6_io_predicateIn_0_valid = Loop_0_io_loopExit_0_valid; // @[bbgemm.scala 331:26]
  assign bb_6_io_predicateIn_0_bits_taskID = Loop_0_io_loopExit_0_bits_taskID; // @[bbgemm.scala 331:26]
  assign bb_6_io_predicateIn_0_bits_control = Loop_0_io_loopExit_0_bits_control; // @[bbgemm.scala 331:26]
  assign bb_6_io_Out_0_ready = const9_io_enable_ready; // @[bbgemm.scala 632:20]
  assign bb_6_io_Out_1_ready = const10_io_enable_ready; // @[bbgemm.scala 634:21]
  assign bb_6_io_Out_2_ready = binaryOp_31_io_enable_ready; // @[bbgemm.scala 636:25]
  assign bb_6_io_Out_3_ready = icmp_32_io_enable_ready; // @[bbgemm.scala 639:21]
  assign bb_6_io_Out_4_ready = br_33_io_enable_ready; // @[bbgemm.scala 642:19]
  assign bb_7_clock = clock;
  assign bb_7_reset = reset;
  assign bb_7_io_predicateIn_0_valid = Loop_1_io_loopExit_0_valid; // @[bbgemm.scala 333:26]
  assign bb_7_io_predicateIn_0_bits_taskID = Loop_1_io_loopExit_0_bits_taskID; // @[bbgemm.scala 333:26]
  assign bb_7_io_predicateIn_0_bits_control = Loop_1_io_loopExit_0_bits_control; // @[bbgemm.scala 333:26]
  assign bb_7_io_Out_0_ready = const11_io_enable_ready; // @[bbgemm.scala 645:21]
  assign bb_7_io_Out_1_ready = const12_io_enable_ready; // @[bbgemm.scala 647:21]
  assign bb_7_io_Out_2_ready = binaryOp_34_io_enable_ready; // @[bbgemm.scala 649:25]
  assign bb_7_io_Out_3_ready = icmp_35_io_enable_ready; // @[bbgemm.scala 652:21]
  assign bb_7_io_Out_4_ready = br_36_io_enable_ready; // @[bbgemm.scala 655:19]
  assign bb_8_clock = clock;
  assign bb_8_reset = reset;
  assign bb_8_io_predicateIn_0_valid = Loop_2_io_loopExit_0_valid; // @[bbgemm.scala 335:26]
  assign bb_8_io_predicateIn_0_bits_taskID = Loop_2_io_loopExit_0_bits_taskID; // @[bbgemm.scala 335:26]
  assign bb_8_io_predicateIn_0_bits_control = Loop_2_io_loopExit_0_bits_control; // @[bbgemm.scala 335:26]
  assign bb_8_io_Out_0_ready = const13_io_enable_ready; // @[bbgemm.scala 658:21]
  assign bb_8_io_Out_1_ready = const14_io_enable_ready; // @[bbgemm.scala 660:21]
  assign bb_8_io_Out_2_ready = binaryOp_37_io_enable_ready; // @[bbgemm.scala 662:25]
  assign bb_8_io_Out_3_ready = icmp_38_io_enable_ready; // @[bbgemm.scala 665:21]
  assign bb_8_io_Out_4_ready = br_39_io_enable_ready; // @[bbgemm.scala 668:19]
  assign bb_9_clock = clock;
  assign bb_9_reset = reset;
  assign bb_9_io_predicateIn_0_valid = Loop_3_io_loopExit_0_valid; // @[bbgemm.scala 337:26]
  assign bb_9_io_predicateIn_0_bits_taskID = Loop_3_io_loopExit_0_bits_taskID; // @[bbgemm.scala 337:26]
  assign bb_9_io_predicateIn_0_bits_control = Loop_3_io_loopExit_0_bits_control; // @[bbgemm.scala 337:26]
  assign bb_9_io_Out_0_ready = const15_io_enable_ready; // @[bbgemm.scala 671:21]
  assign bb_9_io_Out_1_ready = const16_io_enable_ready; // @[bbgemm.scala 673:21]
  assign bb_9_io_Out_2_ready = binaryOp_40_io_enable_ready; // @[bbgemm.scala 675:25]
  assign bb_9_io_Out_3_ready = icmp_41_io_enable_ready; // @[bbgemm.scala 678:21]
  assign bb_9_io_Out_4_ready = br_42_io_enable_ready; // @[bbgemm.scala 681:19]
  assign bb_10_clock = clock;
  assign bb_10_reset = reset;
  assign bb_10_io_predicateIn_0_valid = Loop_4_io_loopExit_0_valid; // @[bbgemm.scala 339:27]
  assign bb_10_io_predicateIn_0_bits_taskID = Loop_4_io_loopExit_0_bits_taskID; // @[bbgemm.scala 339:27]
  assign bb_10_io_predicateIn_0_bits_control = Loop_4_io_loopExit_0_bits_control; // @[bbgemm.scala 339:27]
  assign bb_10_io_Out_0_ready = ret_43_io_In_enable_ready; // @[bbgemm.scala 684:23]
  assign br_0_clock = clock;
  assign br_0_reset = reset;
  assign br_0_io_enable_valid = bb_0_io_Out_0_valid; // @[bbgemm.scala 521:18]
  assign br_0_io_enable_bits_taskID = bb_0_io_Out_0_bits_taskID; // @[bbgemm.scala 521:18]
  assign br_0_io_enable_bits_control = bb_0_io_Out_0_bits_control; // @[bbgemm.scala 521:18]
  assign br_0_io_Out_0_ready = Loop_4_io_enable_ready; // @[bbgemm.scala 377:20]
  assign phi1_clock = clock;
  assign phi1_reset = reset;
  assign phi1_io_enable_valid = bb_1_io_Out_1_valid; // @[bbgemm.scala 526:18]
  assign phi1_io_enable_bits_taskID = bb_1_io_Out_1_bits_taskID; // @[bbgemm.scala 526:18]
  assign phi1_io_enable_bits_control = bb_1_io_Out_1_bits_control; // @[bbgemm.scala 526:18]
  assign phi1_io_InData_0_valid = const0_io_Out_valid; // @[bbgemm.scala 743:21]
  assign phi1_io_InData_0_bits_taskID = const0_io_Out_bits_taskID; // @[bbgemm.scala 743:21]
  assign phi1_io_InData_1_valid = Loop_4_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 513:21]
  assign phi1_io_InData_1_bits_taskID = Loop_4_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 513:21]
  assign phi1_io_InData_1_bits_data = Loop_4_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 513:21]
  assign phi1_io_Mask_valid = bb_1_io_MaskBB_0_valid; // @[bbgemm.scala 693:16]
  assign phi1_io_Mask_bits = bb_1_io_MaskBB_0_bits; // @[bbgemm.scala 693:16]
  assign phi1_io_Out_0_ready = Loop_3_io_InLiveIn_0_ready; // @[bbgemm.scala 429:25]
  assign phi1_io_Out_1_ready = binaryOp_40_io_LeftIO_ready; // @[bbgemm.scala 777:25]
  assign br_2_clock = clock;
  assign br_2_reset = reset;
  assign br_2_io_enable_valid = bb_1_io_Out_2_valid; // @[bbgemm.scala 529:18]
  assign br_2_io_enable_bits_taskID = bb_1_io_Out_2_bits_taskID; // @[bbgemm.scala 529:18]
  assign br_2_io_enable_bits_control = bb_1_io_Out_2_bits_control; // @[bbgemm.scala 529:18]
  assign br_2_io_Out_0_ready = Loop_3_io_enable_ready; // @[bbgemm.scala 371:20]
  assign phi3_clock = clock;
  assign phi3_reset = reset;
  assign phi3_io_enable_valid = bb_2_io_Out_1_valid; // @[bbgemm.scala 534:18]
  assign phi3_io_enable_bits_taskID = bb_2_io_Out_1_bits_taskID; // @[bbgemm.scala 534:18]
  assign phi3_io_enable_bits_control = bb_2_io_Out_1_bits_control; // @[bbgemm.scala 534:18]
  assign phi3_io_InData_0_valid = const1_io_Out_valid; // @[bbgemm.scala 745:21]
  assign phi3_io_InData_0_bits_taskID = const1_io_Out_bits_taskID; // @[bbgemm.scala 745:21]
  assign phi3_io_InData_1_valid = Loop_3_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 511:21]
  assign phi3_io_InData_1_bits_taskID = Loop_3_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 511:21]
  assign phi3_io_InData_1_bits_data = Loop_3_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 511:21]
  assign phi3_io_Mask_valid = bb_2_io_MaskBB_0_valid; // @[bbgemm.scala 695:16]
  assign phi3_io_Mask_bits = bb_2_io_MaskBB_0_bits; // @[bbgemm.scala 695:16]
  assign phi3_io_Out_0_ready = Loop_2_io_InLiveIn_0_ready; // @[bbgemm.scala 419:25]
  assign phi3_io_Out_1_ready = binaryOp_37_io_LeftIO_ready; // @[bbgemm.scala 779:25]
  assign br_4_clock = clock;
  assign br_4_reset = reset;
  assign br_4_io_enable_valid = bb_2_io_Out_2_valid; // @[bbgemm.scala 537:18]
  assign br_4_io_enable_bits_taskID = bb_2_io_Out_2_bits_taskID; // @[bbgemm.scala 537:18]
  assign br_4_io_enable_bits_control = bb_2_io_Out_2_bits_control; // @[bbgemm.scala 537:18]
  assign br_4_io_Out_0_ready = Loop_2_io_enable_ready; // @[bbgemm.scala 365:20]
  assign phi5_clock = clock;
  assign phi5_reset = reset;
  assign phi5_io_enable_valid = bb_3_io_Out_2_valid; // @[bbgemm.scala 544:18]
  assign phi5_io_enable_bits_taskID = bb_3_io_Out_2_bits_taskID; // @[bbgemm.scala 544:18]
  assign phi5_io_enable_bits_control = bb_3_io_Out_2_bits_control; // @[bbgemm.scala 544:18]
  assign phi5_io_InData_0_valid = const2_io_Out_valid; // @[bbgemm.scala 747:21]
  assign phi5_io_InData_0_bits_taskID = const2_io_Out_bits_taskID; // @[bbgemm.scala 747:21]
  assign phi5_io_InData_1_valid = Loop_2_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 509:21]
  assign phi5_io_InData_1_bits_taskID = Loop_2_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 509:21]
  assign phi5_io_InData_1_bits_data = Loop_2_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 509:21]
  assign phi5_io_Mask_valid = bb_3_io_MaskBB_0_valid; // @[bbgemm.scala 697:16]
  assign phi5_io_Mask_bits = bb_3_io_MaskBB_0_bits; // @[bbgemm.scala 697:16]
  assign phi5_io_Out_0_ready = binaryOp_6_io_LeftIO_ready; // @[bbgemm.scala 781:24]
  assign phi5_io_Out_1_ready = binaryOp_34_io_LeftIO_ready; // @[bbgemm.scala 783:25]
  assign binaryOp_6_clock = clock;
  assign binaryOp_6_reset = reset;
  assign binaryOp_6_io_enable_valid = bb_3_io_Out_3_valid; // @[bbgemm.scala 547:24]
  assign binaryOp_6_io_enable_bits_control = bb_3_io_Out_3_bits_control; // @[bbgemm.scala 547:24]
  assign binaryOp_6_io_Out_0_ready = Loop_1_io_InLiveIn_0_ready; // @[bbgemm.scala 407:25]
  assign binaryOp_6_io_LeftIO_valid = phi5_io_Out_0_valid; // @[bbgemm.scala 781:24]
  assign binaryOp_6_io_LeftIO_bits_data = phi5_io_Out_0_bits_data; // @[bbgemm.scala 781:24]
  assign binaryOp_6_io_RightIO_valid = const3_io_Out_valid; // @[bbgemm.scala 749:25]
  assign br_7_clock = clock;
  assign br_7_reset = reset;
  assign br_7_io_enable_valid = bb_3_io_Out_4_valid; // @[bbgemm.scala 550:18]
  assign br_7_io_enable_bits_taskID = bb_3_io_Out_4_bits_taskID; // @[bbgemm.scala 550:18]
  assign br_7_io_enable_bits_control = bb_3_io_Out_4_bits_control; // @[bbgemm.scala 550:18]
  assign br_7_io_Out_0_ready = Loop_1_io_enable_ready; // @[bbgemm.scala 359:20]
  assign phi8_clock = clock;
  assign phi8_reset = reset;
  assign phi8_io_enable_valid = bb_4_io_Out_2_valid; // @[bbgemm.scala 557:18]
  assign phi8_io_enable_bits_taskID = bb_4_io_Out_2_bits_taskID; // @[bbgemm.scala 557:18]
  assign phi8_io_enable_bits_control = bb_4_io_Out_2_bits_control; // @[bbgemm.scala 557:18]
  assign phi8_io_InData_0_valid = const4_io_Out_valid; // @[bbgemm.scala 751:21]
  assign phi8_io_InData_0_bits_taskID = const4_io_Out_bits_taskID; // @[bbgemm.scala 751:21]
  assign phi8_io_InData_1_valid = Loop_1_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 507:21]
  assign phi8_io_InData_1_bits_taskID = Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 507:21]
  assign phi8_io_InData_1_bits_data = Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 507:21]
  assign phi8_io_Mask_valid = bb_4_io_MaskBB_0_valid; // @[bbgemm.scala 699:16]
  assign phi8_io_Mask_bits = bb_4_io_MaskBB_0_bits; // @[bbgemm.scala 699:16]
  assign phi8_io_Out_0_ready = binaryOp_9_io_LeftIO_ready; // @[bbgemm.scala 785:24]
  assign phi8_io_Out_1_ready = binaryOp_11_io_LeftIO_ready; // @[bbgemm.scala 787:25]
  assign phi8_io_Out_2_ready = binaryOp_31_io_LeftIO_ready; // @[bbgemm.scala 789:25]
  assign binaryOp_9_clock = clock;
  assign binaryOp_9_reset = reset;
  assign binaryOp_9_io_enable_valid = bb_4_io_Out_3_valid; // @[bbgemm.scala 560:24]
  assign binaryOp_9_io_enable_bits_control = bb_4_io_Out_3_bits_control; // @[bbgemm.scala 560:24]
  assign binaryOp_9_io_Out_0_ready = binaryOp_10_io_LeftIO_ready; // @[bbgemm.scala 791:25]
  assign binaryOp_9_io_LeftIO_valid = phi8_io_Out_0_valid; // @[bbgemm.scala 785:24]
  assign binaryOp_9_io_LeftIO_bits_data = phi8_io_Out_0_bits_data; // @[bbgemm.scala 785:24]
  assign binaryOp_9_io_RightIO_valid = Loop_1_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 465:25]
  assign binaryOp_9_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 465:25]
  assign binaryOp_10_clock = clock;
  assign binaryOp_10_reset = reset;
  assign binaryOp_10_io_enable_valid = bb_4_io_Out_4_valid; // @[bbgemm.scala 563:25]
  assign binaryOp_10_io_enable_bits_control = bb_4_io_Out_4_bits_control; // @[bbgemm.scala 563:25]
  assign binaryOp_10_io_Out_0_ready = Loop_0_io_InLiveIn_0_ready; // @[bbgemm.scala 395:25]
  assign binaryOp_10_io_LeftIO_valid = binaryOp_9_io_Out_0_valid; // @[bbgemm.scala 791:25]
  assign binaryOp_10_io_LeftIO_bits_data = binaryOp_9_io_Out_0_bits_data; // @[bbgemm.scala 791:25]
  assign binaryOp_10_io_RightIO_valid = const5_io_Out_valid; // @[bbgemm.scala 753:26]
  assign binaryOp_11_clock = clock;
  assign binaryOp_11_reset = reset;
  assign binaryOp_11_io_enable_valid = bb_4_io_Out_5_valid; // @[bbgemm.scala 566:25]
  assign binaryOp_11_io_enable_bits_control = bb_4_io_Out_5_bits_control; // @[bbgemm.scala 566:25]
  assign binaryOp_11_io_Out_0_ready = binaryOp_12_io_LeftIO_ready; // @[bbgemm.scala 793:25]
  assign binaryOp_11_io_LeftIO_valid = phi8_io_Out_1_valid; // @[bbgemm.scala 787:25]
  assign binaryOp_11_io_LeftIO_bits_data = phi8_io_Out_1_bits_data; // @[bbgemm.scala 787:25]
  assign binaryOp_11_io_RightIO_valid = Loop_1_io_OutLiveIn_field4_1_valid; // @[bbgemm.scala 467:26]
  assign binaryOp_11_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field4_1_bits_data; // @[bbgemm.scala 467:26]
  assign binaryOp_12_clock = clock;
  assign binaryOp_12_reset = reset;
  assign binaryOp_12_io_enable_valid = bb_4_io_Out_6_valid; // @[bbgemm.scala 569:25]
  assign binaryOp_12_io_enable_bits_control = bb_4_io_Out_6_bits_control; // @[bbgemm.scala 569:25]
  assign binaryOp_12_io_Out_0_ready = Gep_13_io_idx_0_ready; // @[bbgemm.scala 795:20]
  assign binaryOp_12_io_LeftIO_valid = binaryOp_11_io_Out_0_valid; // @[bbgemm.scala 793:25]
  assign binaryOp_12_io_LeftIO_bits_data = binaryOp_11_io_Out_0_bits_data; // @[bbgemm.scala 793:25]
  assign binaryOp_12_io_RightIO_valid = Loop_1_io_OutLiveIn_field0_1_valid; // @[bbgemm.scala 463:26]
  assign binaryOp_12_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field0_1_bits_data; // @[bbgemm.scala 463:26]
  assign Gep_13_clock = clock;
  assign Gep_13_reset = reset;
  assign Gep_13_io_enable_valid = bb_4_io_Out_7_valid; // @[bbgemm.scala 572:20]
  assign Gep_13_io_enable_bits_control = bb_4_io_Out_7_bits_control; // @[bbgemm.scala 572:20]
  assign Gep_13_io_Out_0_ready = ld_14_io_GepAddr_ready; // @[bbgemm.scala 797:20]
  assign Gep_13_io_baseAddress_valid = Loop_1_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 469:25]
  assign Gep_13_io_baseAddress_bits_taskID = Loop_1_io_OutLiveIn_field5_0_bits_taskID; // @[bbgemm.scala 469:25]
  assign Gep_13_io_baseAddress_bits_data = Loop_1_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 469:25]
  assign Gep_13_io_idx_0_valid = binaryOp_12_io_Out_0_valid; // @[bbgemm.scala 795:20]
  assign Gep_13_io_idx_0_bits_data = binaryOp_12_io_Out_0_bits_data; // @[bbgemm.scala 795:20]
  assign ld_14_clock = clock;
  assign ld_14_reset = reset;
  assign ld_14_io_enable_valid = bb_4_io_Out_8_valid; // @[bbgemm.scala 575:19]
  assign ld_14_io_enable_bits_taskID = bb_4_io_Out_8_bits_taskID; // @[bbgemm.scala 575:19]
  assign ld_14_io_enable_bits_control = bb_4_io_Out_8_bits_control; // @[bbgemm.scala 575:19]
  assign ld_14_io_Out_0_ready = Loop_0_io_InLiveIn_1_ready; // @[bbgemm.scala 397:25]
  assign ld_14_io_GepAddr_valid = Gep_13_io_Out_0_valid; // @[bbgemm.scala 797:20]
  assign ld_14_io_GepAddr_bits_predicate = Gep_13_io_Out_0_bits_predicate; // @[bbgemm.scala 797:20]
  assign ld_14_io_GepAddr_bits_taskID = Gep_13_io_Out_0_bits_taskID; // @[bbgemm.scala 797:20]
  assign ld_14_io_GepAddr_bits_data = Gep_13_io_Out_0_bits_data; // @[bbgemm.scala 797:20]
  assign ld_14_io_memReq_ready = MemCtrl_io_ReadIn_0_ready; // @[bbgemm.scala 715:24]
  assign ld_14_io_memResp_valid = MemCtrl_io_ReadOut_0_valid; // @[bbgemm.scala 717:20]
  assign ld_14_io_memResp_data = MemCtrl_io_ReadOut_0_data; // @[bbgemm.scala 717:20]
  assign br_15_clock = clock;
  assign br_15_reset = reset;
  assign br_15_io_enable_valid = bb_4_io_Out_9_valid; // @[bbgemm.scala 578:19]
  assign br_15_io_enable_bits_taskID = bb_4_io_Out_9_bits_taskID; // @[bbgemm.scala 578:19]
  assign br_15_io_enable_bits_control = bb_4_io_Out_9_bits_control; // @[bbgemm.scala 578:19]
  assign br_15_io_Out_0_ready = Loop_0_io_enable_ready; // @[bbgemm.scala 353:20]
  assign phi16_clock = clock;
  assign phi16_reset = reset;
  assign phi16_io_enable_valid = bb_5_io_Out_3_valid; // @[bbgemm.scala 587:19]
  assign phi16_io_enable_bits_taskID = bb_5_io_Out_3_bits_taskID; // @[bbgemm.scala 587:19]
  assign phi16_io_enable_bits_control = bb_5_io_Out_3_bits_control; // @[bbgemm.scala 587:19]
  assign phi16_io_InData_0_valid = const6_io_Out_valid; // @[bbgemm.scala 755:22]
  assign phi16_io_InData_0_bits_taskID = const6_io_Out_bits_taskID; // @[bbgemm.scala 755:22]
  assign phi16_io_InData_1_valid = Loop_0_io_CarryDepenOut_field0_0_valid; // @[bbgemm.scala 505:22]
  assign phi16_io_InData_1_bits_taskID = Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[bbgemm.scala 505:22]
  assign phi16_io_InData_1_bits_data = Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[bbgemm.scala 505:22]
  assign phi16_io_Mask_valid = bb_5_io_MaskBB_0_valid; // @[bbgemm.scala 701:17]
  assign phi16_io_Mask_bits = bb_5_io_MaskBB_0_bits; // @[bbgemm.scala 701:17]
  assign phi16_io_Out_0_ready = binaryOp_17_io_LeftIO_ready; // @[bbgemm.scala 799:25]
  assign phi16_io_Out_1_ready = binaryOp_22_io_LeftIO_ready; // @[bbgemm.scala 801:25]
  assign phi16_io_Out_2_ready = binaryOp_28_io_LeftIO_ready; // @[bbgemm.scala 803:25]
  assign binaryOp_17_clock = clock;
  assign binaryOp_17_reset = reset;
  assign binaryOp_17_io_enable_valid = bb_5_io_Out_4_valid; // @[bbgemm.scala 590:25]
  assign binaryOp_17_io_enable_bits_control = bb_5_io_Out_4_bits_control; // @[bbgemm.scala 590:25]
  assign binaryOp_17_io_Out_0_ready = binaryOp_18_io_LeftIO_ready; // @[bbgemm.scala 805:25]
  assign binaryOp_17_io_LeftIO_valid = phi16_io_Out_0_valid; // @[bbgemm.scala 799:25]
  assign binaryOp_17_io_LeftIO_bits_data = phi16_io_Out_0_bits_data; // @[bbgemm.scala 799:25]
  assign binaryOp_17_io_RightIO_valid = Loop_0_io_OutLiveIn_field5_0_valid; // @[bbgemm.scala 459:26]
  assign binaryOp_17_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field5_0_bits_data; // @[bbgemm.scala 459:26]
  assign binaryOp_18_clock = clock;
  assign binaryOp_18_reset = reset;
  assign binaryOp_18_io_enable_valid = bb_5_io_Out_5_valid; // @[bbgemm.scala 593:25]
  assign binaryOp_18_io_enable_bits_control = bb_5_io_Out_5_bits_control; // @[bbgemm.scala 593:25]
  assign binaryOp_18_io_Out_0_ready = Gep_19_io_idx_0_ready; // @[bbgemm.scala 807:20]
  assign binaryOp_18_io_LeftIO_valid = binaryOp_17_io_Out_0_valid; // @[bbgemm.scala 805:25]
  assign binaryOp_18_io_LeftIO_bits_data = binaryOp_17_io_Out_0_bits_data; // @[bbgemm.scala 805:25]
  assign binaryOp_18_io_RightIO_valid = Loop_0_io_OutLiveIn_field0_0_valid; // @[bbgemm.scala 449:26]
  assign binaryOp_18_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field0_0_bits_data; // @[bbgemm.scala 449:26]
  assign Gep_19_clock = clock;
  assign Gep_19_reset = reset;
  assign Gep_19_io_enable_valid = bb_5_io_Out_6_valid; // @[bbgemm.scala 596:20]
  assign Gep_19_io_enable_bits_control = bb_5_io_Out_6_bits_control; // @[bbgemm.scala 596:20]
  assign Gep_19_io_Out_0_ready = ld_20_io_GepAddr_ready; // @[bbgemm.scala 809:20]
  assign Gep_19_io_baseAddress_valid = Loop_0_io_OutLiveIn_field4_0_valid; // @[bbgemm.scala 457:25]
  assign Gep_19_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field4_0_bits_taskID; // @[bbgemm.scala 457:25]
  assign Gep_19_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field4_0_bits_data; // @[bbgemm.scala 457:25]
  assign Gep_19_io_idx_0_valid = binaryOp_18_io_Out_0_valid; // @[bbgemm.scala 807:20]
  assign Gep_19_io_idx_0_bits_data = binaryOp_18_io_Out_0_bits_data; // @[bbgemm.scala 807:20]
  assign ld_20_clock = clock;
  assign ld_20_reset = reset;
  assign ld_20_io_enable_valid = bb_5_io_Out_7_valid; // @[bbgemm.scala 599:19]
  assign ld_20_io_enable_bits_taskID = bb_5_io_Out_7_bits_taskID; // @[bbgemm.scala 599:19]
  assign ld_20_io_enable_bits_control = bb_5_io_Out_7_bits_control; // @[bbgemm.scala 599:19]
  assign ld_20_io_Out_0_ready = FP_21_io_RightIO_ready; // @[bbgemm.scala 811:20]
  assign ld_20_io_GepAddr_valid = Gep_19_io_Out_0_valid; // @[bbgemm.scala 809:20]
  assign ld_20_io_GepAddr_bits_predicate = Gep_19_io_Out_0_bits_predicate; // @[bbgemm.scala 809:20]
  assign ld_20_io_GepAddr_bits_taskID = Gep_19_io_Out_0_bits_taskID; // @[bbgemm.scala 809:20]
  assign ld_20_io_GepAddr_bits_data = Gep_19_io_Out_0_bits_data; // @[bbgemm.scala 809:20]
  assign ld_20_io_memReq_ready = MemCtrl_io_ReadIn_1_ready; // @[bbgemm.scala 719:24]
  assign ld_20_io_memResp_valid = MemCtrl_io_ReadOut_1_valid; // @[bbgemm.scala 721:20]
  assign ld_20_io_memResp_data = MemCtrl_io_ReadOut_1_data; // @[bbgemm.scala 721:20]
  assign FP_21_clock = clock;
  assign FP_21_reset = reset;
  assign FP_21_io_enable_valid = bb_5_io_Out_8_valid; // @[bbgemm.scala 602:19]
  assign FP_21_io_enable_bits_taskID = bb_5_io_Out_8_bits_taskID; // @[bbgemm.scala 602:19]
  assign FP_21_io_enable_bits_control = bb_5_io_Out_8_bits_control; // @[bbgemm.scala 602:19]
  assign FP_21_io_Out_0_ready = FP_26_io_RightIO_ready; // @[bbgemm.scala 813:20]
  assign FP_21_io_LeftIO_valid = Loop_0_io_OutLiveIn_field1_0_valid; // @[bbgemm.scala 451:19]
  assign FP_21_io_LeftIO_bits_taskID = Loop_0_io_OutLiveIn_field1_0_bits_taskID; // @[bbgemm.scala 451:19]
  assign FP_21_io_LeftIO_bits_data = Loop_0_io_OutLiveIn_field1_0_bits_data; // @[bbgemm.scala 451:19]
  assign FP_21_io_RightIO_valid = ld_20_io_Out_0_valid; // @[bbgemm.scala 811:20]
  assign FP_21_io_RightIO_bits_taskID = ld_20_io_Out_0_bits_taskID; // @[bbgemm.scala 811:20]
  assign FP_21_io_RightIO_bits_data = ld_20_io_Out_0_bits_data; // @[bbgemm.scala 811:20]
  assign binaryOp_22_clock = clock;
  assign binaryOp_22_reset = reset;
  assign binaryOp_22_io_enable_valid = bb_5_io_Out_9_valid; // @[bbgemm.scala 605:25]
  assign binaryOp_22_io_enable_bits_control = bb_5_io_Out_9_bits_control; // @[bbgemm.scala 605:25]
  assign binaryOp_22_io_Out_0_ready = binaryOp_23_io_LeftIO_ready; // @[bbgemm.scala 815:25]
  assign binaryOp_22_io_LeftIO_valid = phi16_io_Out_1_valid; // @[bbgemm.scala 801:25]
  assign binaryOp_22_io_LeftIO_bits_data = phi16_io_Out_1_bits_data; // @[bbgemm.scala 801:25]
  assign binaryOp_22_io_RightIO_valid = Loop_0_io_OutLiveIn_field5_1_valid; // @[bbgemm.scala 461:26]
  assign binaryOp_22_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field5_1_bits_data; // @[bbgemm.scala 461:26]
  assign binaryOp_23_clock = clock;
  assign binaryOp_23_reset = reset;
  assign binaryOp_23_io_enable_valid = bb_5_io_Out_10_valid; // @[bbgemm.scala 608:25]
  assign binaryOp_23_io_enable_bits_control = bb_5_io_Out_10_bits_control; // @[bbgemm.scala 608:25]
  assign binaryOp_23_io_Out_0_ready = Gep_24_io_idx_0_ready; // @[bbgemm.scala 817:20]
  assign binaryOp_23_io_LeftIO_valid = binaryOp_22_io_Out_0_valid; // @[bbgemm.scala 815:25]
  assign binaryOp_23_io_LeftIO_bits_data = binaryOp_22_io_Out_0_bits_data; // @[bbgemm.scala 815:25]
  assign binaryOp_23_io_RightIO_valid = Loop_0_io_OutLiveIn_field2_0_valid; // @[bbgemm.scala 453:26]
  assign binaryOp_23_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field2_0_bits_data; // @[bbgemm.scala 453:26]
  assign Gep_24_clock = clock;
  assign Gep_24_reset = reset;
  assign Gep_24_io_enable_valid = bb_5_io_Out_11_valid; // @[bbgemm.scala 611:20]
  assign Gep_24_io_enable_bits_control = bb_5_io_Out_11_bits_control; // @[bbgemm.scala 611:20]
  assign Gep_24_io_Out_0_ready = ld_25_io_GepAddr_ready; // @[bbgemm.scala 819:20]
  assign Gep_24_io_Out_1_ready = st_27_io_GepAddr_ready; // @[bbgemm.scala 821:20]
  assign Gep_24_io_baseAddress_valid = Loop_0_io_OutLiveIn_field3_0_valid; // @[bbgemm.scala 455:25]
  assign Gep_24_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field3_0_bits_taskID; // @[bbgemm.scala 455:25]
  assign Gep_24_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field3_0_bits_data; // @[bbgemm.scala 455:25]
  assign Gep_24_io_idx_0_valid = binaryOp_23_io_Out_0_valid; // @[bbgemm.scala 817:20]
  assign Gep_24_io_idx_0_bits_data = binaryOp_23_io_Out_0_bits_data; // @[bbgemm.scala 817:20]
  assign ld_25_clock = clock;
  assign ld_25_reset = reset;
  assign ld_25_io_enable_valid = bb_5_io_Out_12_valid; // @[bbgemm.scala 614:19]
  assign ld_25_io_enable_bits_taskID = bb_5_io_Out_12_bits_taskID; // @[bbgemm.scala 614:19]
  assign ld_25_io_enable_bits_control = bb_5_io_Out_12_bits_control; // @[bbgemm.scala 614:19]
  assign ld_25_io_Out_0_ready = FP_26_io_LeftIO_ready; // @[bbgemm.scala 823:19]
  assign ld_25_io_GepAddr_valid = Gep_24_io_Out_0_valid; // @[bbgemm.scala 819:20]
  assign ld_25_io_GepAddr_bits_predicate = Gep_24_io_Out_0_bits_predicate; // @[bbgemm.scala 819:20]
  assign ld_25_io_GepAddr_bits_taskID = Gep_24_io_Out_0_bits_taskID; // @[bbgemm.scala 819:20]
  assign ld_25_io_GepAddr_bits_data = Gep_24_io_Out_0_bits_data; // @[bbgemm.scala 819:20]
  assign ld_25_io_memReq_ready = MemCtrl_io_ReadIn_2_ready; // @[bbgemm.scala 723:24]
  assign ld_25_io_memResp_valid = MemCtrl_io_ReadOut_2_valid; // @[bbgemm.scala 725:20]
  assign ld_25_io_memResp_data = MemCtrl_io_ReadOut_2_data; // @[bbgemm.scala 725:20]
  assign FP_26_clock = clock;
  assign FP_26_reset = reset;
  assign FP_26_io_enable_valid = bb_5_io_Out_13_valid; // @[bbgemm.scala 617:19]
  assign FP_26_io_enable_bits_taskID = bb_5_io_Out_13_bits_taskID; // @[bbgemm.scala 617:19]
  assign FP_26_io_enable_bits_control = bb_5_io_Out_13_bits_control; // @[bbgemm.scala 617:19]
  assign FP_26_io_Out_0_ready = st_27_io_inData_ready; // @[bbgemm.scala 825:19]
  assign FP_26_io_LeftIO_valid = ld_25_io_Out_0_valid; // @[bbgemm.scala 823:19]
  assign FP_26_io_LeftIO_bits_taskID = ld_25_io_Out_0_bits_taskID; // @[bbgemm.scala 823:19]
  assign FP_26_io_LeftIO_bits_data = ld_25_io_Out_0_bits_data; // @[bbgemm.scala 823:19]
  assign FP_26_io_RightIO_valid = FP_21_io_Out_0_valid; // @[bbgemm.scala 813:20]
  assign FP_26_io_RightIO_bits_taskID = FP_21_io_Out_0_bits_taskID; // @[bbgemm.scala 813:20]
  assign FP_26_io_RightIO_bits_data = FP_21_io_Out_0_bits_data; // @[bbgemm.scala 813:20]
  assign st_27_clock = clock;
  assign st_27_reset = reset;
  assign st_27_io_enable_valid = bb_5_io_Out_14_valid; // @[bbgemm.scala 620:19]
  assign st_27_io_enable_bits_taskID = bb_5_io_Out_14_bits_taskID; // @[bbgemm.scala 620:19]
  assign st_27_io_enable_bits_control = bb_5_io_Out_14_bits_control; // @[bbgemm.scala 620:19]
  assign st_27_io_GepAddr_valid = Gep_24_io_Out_1_valid; // @[bbgemm.scala 821:20]
  assign st_27_io_GepAddr_bits_taskID = Gep_24_io_Out_1_bits_taskID; // @[bbgemm.scala 821:20]
  assign st_27_io_GepAddr_bits_data = Gep_24_io_Out_1_bits_data; // @[bbgemm.scala 821:20]
  assign st_27_io_inData_valid = FP_26_io_Out_0_valid; // @[bbgemm.scala 825:19]
  assign st_27_io_inData_bits_taskID = FP_26_io_Out_0_bits_taskID; // @[bbgemm.scala 825:19]
  assign st_27_io_inData_bits_data = FP_26_io_Out_0_bits_data; // @[bbgemm.scala 825:19]
  assign st_27_io_memReq_ready = MemCtrl_io_WriteIn_0_ready; // @[bbgemm.scala 727:25]
  assign st_27_io_memResp_valid = MemCtrl_io_WriteOut_0_valid; // @[bbgemm.scala 729:20]
  assign binaryOp_28_clock = clock;
  assign binaryOp_28_reset = reset;
  assign binaryOp_28_io_enable_valid = bb_5_io_Out_15_valid; // @[bbgemm.scala 623:25]
  assign binaryOp_28_io_enable_bits_taskID = bb_5_io_Out_15_bits_taskID; // @[bbgemm.scala 623:25]
  assign binaryOp_28_io_enable_bits_control = bb_5_io_Out_15_bits_control; // @[bbgemm.scala 623:25]
  assign binaryOp_28_io_Out_0_ready = Loop_0_io_CarryDepenIn_0_ready; // @[bbgemm.scala 489:29]
  assign binaryOp_28_io_Out_1_ready = icmp_29_io_LeftIO_ready; // @[bbgemm.scala 827:21]
  assign binaryOp_28_io_LeftIO_valid = phi16_io_Out_2_valid; // @[bbgemm.scala 803:25]
  assign binaryOp_28_io_LeftIO_bits_taskID = phi16_io_Out_2_bits_taskID; // @[bbgemm.scala 803:25]
  assign binaryOp_28_io_LeftIO_bits_data = phi16_io_Out_2_bits_data; // @[bbgemm.scala 803:25]
  assign binaryOp_28_io_RightIO_valid = const7_io_Out_valid; // @[bbgemm.scala 757:26]
  assign binaryOp_28_io_RightIO_bits_taskID = const7_io_Out_bits_taskID; // @[bbgemm.scala 757:26]
  assign icmp_29_clock = clock;
  assign icmp_29_reset = reset;
  assign icmp_29_io_enable_valid = bb_5_io_Out_16_valid; // @[bbgemm.scala 626:21]
  assign icmp_29_io_enable_bits_taskID = bb_5_io_Out_16_bits_taskID; // @[bbgemm.scala 626:21]
  assign icmp_29_io_enable_bits_control = bb_5_io_Out_16_bits_control; // @[bbgemm.scala 626:21]
  assign icmp_29_io_Out_0_ready = br_30_io_CmpIO_ready; // @[bbgemm.scala 829:18]
  assign icmp_29_io_LeftIO_valid = binaryOp_28_io_Out_1_valid; // @[bbgemm.scala 827:21]
  assign icmp_29_io_LeftIO_bits_taskID = binaryOp_28_io_Out_1_bits_taskID; // @[bbgemm.scala 827:21]
  assign icmp_29_io_LeftIO_bits_data = binaryOp_28_io_Out_1_bits_data; // @[bbgemm.scala 827:21]
  assign icmp_29_io_RightIO_valid = const8_io_Out_valid; // @[bbgemm.scala 759:22]
  assign icmp_29_io_RightIO_bits_taskID = const8_io_Out_bits_taskID; // @[bbgemm.scala 759:22]
  assign br_30_clock = clock;
  assign br_30_reset = reset;
  assign br_30_io_enable_valid = bb_5_io_Out_17_valid; // @[bbgemm.scala 629:19]
  assign br_30_io_enable_bits_taskID = bb_5_io_Out_17_bits_taskID; // @[bbgemm.scala 629:19]
  assign br_30_io_enable_bits_control = bb_5_io_Out_17_bits_control; // @[bbgemm.scala 629:19]
  assign br_30_io_CmpIO_valid = icmp_29_io_Out_0_valid; // @[bbgemm.scala 829:18]
  assign br_30_io_CmpIO_bits_taskID = icmp_29_io_Out_0_bits_taskID; // @[bbgemm.scala 829:18]
  assign br_30_io_CmpIO_bits_data = icmp_29_io_Out_0_bits_data; // @[bbgemm.scala 829:18]
  assign br_30_io_TrueOutput_0_ready = Loop_0_io_loopFinish_0_ready; // @[bbgemm.scala 357:27]
  assign br_30_io_FalseOutput_0_ready = Loop_0_io_loopBack_0_ready; // @[bbgemm.scala 355:25]
  assign binaryOp_31_clock = clock;
  assign binaryOp_31_reset = reset;
  assign binaryOp_31_io_enable_valid = bb_6_io_Out_2_valid; // @[bbgemm.scala 636:25]
  assign binaryOp_31_io_enable_bits_taskID = bb_6_io_Out_2_bits_taskID; // @[bbgemm.scala 636:25]
  assign binaryOp_31_io_enable_bits_control = bb_6_io_Out_2_bits_control; // @[bbgemm.scala 636:25]
  assign binaryOp_31_io_Out_0_ready = Loop_1_io_CarryDepenIn_0_ready; // @[bbgemm.scala 491:29]
  assign binaryOp_31_io_Out_1_ready = icmp_32_io_LeftIO_ready; // @[bbgemm.scala 831:21]
  assign binaryOp_31_io_LeftIO_valid = phi8_io_Out_2_valid; // @[bbgemm.scala 789:25]
  assign binaryOp_31_io_LeftIO_bits_taskID = phi8_io_Out_2_bits_taskID; // @[bbgemm.scala 789:25]
  assign binaryOp_31_io_LeftIO_bits_data = phi8_io_Out_2_bits_data; // @[bbgemm.scala 789:25]
  assign binaryOp_31_io_RightIO_valid = const9_io_Out_valid; // @[bbgemm.scala 761:26]
  assign binaryOp_31_io_RightIO_bits_taskID = const9_io_Out_bits_taskID; // @[bbgemm.scala 761:26]
  assign icmp_32_clock = clock;
  assign icmp_32_reset = reset;
  assign icmp_32_io_enable_valid = bb_6_io_Out_3_valid; // @[bbgemm.scala 639:21]
  assign icmp_32_io_enable_bits_taskID = bb_6_io_Out_3_bits_taskID; // @[bbgemm.scala 639:21]
  assign icmp_32_io_enable_bits_control = bb_6_io_Out_3_bits_control; // @[bbgemm.scala 639:21]
  assign icmp_32_io_Out_0_ready = br_33_io_CmpIO_ready; // @[bbgemm.scala 833:18]
  assign icmp_32_io_LeftIO_valid = binaryOp_31_io_Out_1_valid; // @[bbgemm.scala 831:21]
  assign icmp_32_io_LeftIO_bits_taskID = binaryOp_31_io_Out_1_bits_taskID; // @[bbgemm.scala 831:21]
  assign icmp_32_io_LeftIO_bits_data = binaryOp_31_io_Out_1_bits_data; // @[bbgemm.scala 831:21]
  assign icmp_32_io_RightIO_valid = const10_io_Out_valid; // @[bbgemm.scala 763:22]
  assign icmp_32_io_RightIO_bits_taskID = const10_io_Out_bits_taskID; // @[bbgemm.scala 763:22]
  assign br_33_clock = clock;
  assign br_33_reset = reset;
  assign br_33_io_enable_valid = bb_6_io_Out_4_valid; // @[bbgemm.scala 642:19]
  assign br_33_io_enable_bits_taskID = bb_6_io_Out_4_bits_taskID; // @[bbgemm.scala 642:19]
  assign br_33_io_enable_bits_control = bb_6_io_Out_4_bits_control; // @[bbgemm.scala 642:19]
  assign br_33_io_CmpIO_valid = icmp_32_io_Out_0_valid; // @[bbgemm.scala 833:18]
  assign br_33_io_CmpIO_bits_taskID = icmp_32_io_Out_0_bits_taskID; // @[bbgemm.scala 833:18]
  assign br_33_io_CmpIO_bits_data = icmp_32_io_Out_0_bits_data; // @[bbgemm.scala 833:18]
  assign br_33_io_TrueOutput_0_ready = Loop_1_io_loopFinish_0_ready; // @[bbgemm.scala 363:27]
  assign br_33_io_FalseOutput_0_ready = Loop_1_io_loopBack_0_ready; // @[bbgemm.scala 361:25]
  assign binaryOp_34_clock = clock;
  assign binaryOp_34_reset = reset;
  assign binaryOp_34_io_enable_valid = bb_7_io_Out_2_valid; // @[bbgemm.scala 649:25]
  assign binaryOp_34_io_enable_bits_taskID = bb_7_io_Out_2_bits_taskID; // @[bbgemm.scala 649:25]
  assign binaryOp_34_io_enable_bits_control = bb_7_io_Out_2_bits_control; // @[bbgemm.scala 649:25]
  assign binaryOp_34_io_Out_0_ready = Loop_2_io_CarryDepenIn_0_ready; // @[bbgemm.scala 493:29]
  assign binaryOp_34_io_Out_1_ready = icmp_35_io_LeftIO_ready; // @[bbgemm.scala 835:21]
  assign binaryOp_34_io_LeftIO_valid = phi5_io_Out_1_valid; // @[bbgemm.scala 783:25]
  assign binaryOp_34_io_LeftIO_bits_taskID = phi5_io_Out_1_bits_taskID; // @[bbgemm.scala 783:25]
  assign binaryOp_34_io_LeftIO_bits_data = phi5_io_Out_1_bits_data; // @[bbgemm.scala 783:25]
  assign binaryOp_34_io_RightIO_valid = const11_io_Out_valid; // @[bbgemm.scala 765:26]
  assign binaryOp_34_io_RightIO_bits_taskID = const11_io_Out_bits_taskID; // @[bbgemm.scala 765:26]
  assign icmp_35_clock = clock;
  assign icmp_35_reset = reset;
  assign icmp_35_io_enable_valid = bb_7_io_Out_3_valid; // @[bbgemm.scala 652:21]
  assign icmp_35_io_enable_bits_taskID = bb_7_io_Out_3_bits_taskID; // @[bbgemm.scala 652:21]
  assign icmp_35_io_enable_bits_control = bb_7_io_Out_3_bits_control; // @[bbgemm.scala 652:21]
  assign icmp_35_io_Out_0_ready = br_36_io_CmpIO_ready; // @[bbgemm.scala 837:18]
  assign icmp_35_io_LeftIO_valid = binaryOp_34_io_Out_1_valid; // @[bbgemm.scala 835:21]
  assign icmp_35_io_LeftIO_bits_taskID = binaryOp_34_io_Out_1_bits_taskID; // @[bbgemm.scala 835:21]
  assign icmp_35_io_LeftIO_bits_data = binaryOp_34_io_Out_1_bits_data; // @[bbgemm.scala 835:21]
  assign icmp_35_io_RightIO_valid = const12_io_Out_valid; // @[bbgemm.scala 767:22]
  assign icmp_35_io_RightIO_bits_taskID = const12_io_Out_bits_taskID; // @[bbgemm.scala 767:22]
  assign br_36_clock = clock;
  assign br_36_reset = reset;
  assign br_36_io_enable_valid = bb_7_io_Out_4_valid; // @[bbgemm.scala 655:19]
  assign br_36_io_enable_bits_taskID = bb_7_io_Out_4_bits_taskID; // @[bbgemm.scala 655:19]
  assign br_36_io_enable_bits_control = bb_7_io_Out_4_bits_control; // @[bbgemm.scala 655:19]
  assign br_36_io_CmpIO_valid = icmp_35_io_Out_0_valid; // @[bbgemm.scala 837:18]
  assign br_36_io_CmpIO_bits_taskID = icmp_35_io_Out_0_bits_taskID; // @[bbgemm.scala 837:18]
  assign br_36_io_CmpIO_bits_data = icmp_35_io_Out_0_bits_data; // @[bbgemm.scala 837:18]
  assign br_36_io_TrueOutput_0_ready = Loop_2_io_loopFinish_0_ready; // @[bbgemm.scala 369:27]
  assign br_36_io_FalseOutput_0_ready = Loop_2_io_loopBack_0_ready; // @[bbgemm.scala 367:25]
  assign binaryOp_37_clock = clock;
  assign binaryOp_37_reset = reset;
  assign binaryOp_37_io_enable_valid = bb_8_io_Out_2_valid; // @[bbgemm.scala 662:25]
  assign binaryOp_37_io_enable_bits_taskID = bb_8_io_Out_2_bits_taskID; // @[bbgemm.scala 662:25]
  assign binaryOp_37_io_enable_bits_control = bb_8_io_Out_2_bits_control; // @[bbgemm.scala 662:25]
  assign binaryOp_37_io_Out_0_ready = Loop_3_io_CarryDepenIn_0_ready; // @[bbgemm.scala 495:29]
  assign binaryOp_37_io_Out_1_ready = icmp_38_io_LeftIO_ready; // @[bbgemm.scala 839:21]
  assign binaryOp_37_io_LeftIO_valid = phi3_io_Out_1_valid; // @[bbgemm.scala 779:25]
  assign binaryOp_37_io_LeftIO_bits_taskID = phi3_io_Out_1_bits_taskID; // @[bbgemm.scala 779:25]
  assign binaryOp_37_io_LeftIO_bits_data = phi3_io_Out_1_bits_data; // @[bbgemm.scala 779:25]
  assign binaryOp_37_io_RightIO_valid = const13_io_Out_valid; // @[bbgemm.scala 769:26]
  assign binaryOp_37_io_RightIO_bits_taskID = const13_io_Out_bits_taskID; // @[bbgemm.scala 769:26]
  assign icmp_38_clock = clock;
  assign icmp_38_reset = reset;
  assign icmp_38_io_enable_valid = bb_8_io_Out_3_valid; // @[bbgemm.scala 665:21]
  assign icmp_38_io_enable_bits_taskID = bb_8_io_Out_3_bits_taskID; // @[bbgemm.scala 665:21]
  assign icmp_38_io_enable_bits_control = bb_8_io_Out_3_bits_control; // @[bbgemm.scala 665:21]
  assign icmp_38_io_Out_0_ready = br_39_io_CmpIO_ready; // @[bbgemm.scala 841:18]
  assign icmp_38_io_LeftIO_valid = binaryOp_37_io_Out_1_valid; // @[bbgemm.scala 839:21]
  assign icmp_38_io_LeftIO_bits_taskID = binaryOp_37_io_Out_1_bits_taskID; // @[bbgemm.scala 839:21]
  assign icmp_38_io_LeftIO_bits_data = binaryOp_37_io_Out_1_bits_data; // @[bbgemm.scala 839:21]
  assign icmp_38_io_RightIO_valid = const14_io_Out_valid; // @[bbgemm.scala 771:22]
  assign icmp_38_io_RightIO_bits_taskID = const14_io_Out_bits_taskID; // @[bbgemm.scala 771:22]
  assign br_39_clock = clock;
  assign br_39_reset = reset;
  assign br_39_io_enable_valid = bb_8_io_Out_4_valid; // @[bbgemm.scala 668:19]
  assign br_39_io_enable_bits_taskID = bb_8_io_Out_4_bits_taskID; // @[bbgemm.scala 668:19]
  assign br_39_io_enable_bits_control = bb_8_io_Out_4_bits_control; // @[bbgemm.scala 668:19]
  assign br_39_io_CmpIO_valid = icmp_38_io_Out_0_valid; // @[bbgemm.scala 841:18]
  assign br_39_io_CmpIO_bits_taskID = icmp_38_io_Out_0_bits_taskID; // @[bbgemm.scala 841:18]
  assign br_39_io_CmpIO_bits_data = icmp_38_io_Out_0_bits_data; // @[bbgemm.scala 841:18]
  assign br_39_io_TrueOutput_0_ready = Loop_3_io_loopBack_0_ready; // @[bbgemm.scala 373:25]
  assign br_39_io_FalseOutput_0_ready = Loop_3_io_loopFinish_0_ready; // @[bbgemm.scala 375:27]
  assign binaryOp_40_clock = clock;
  assign binaryOp_40_reset = reset;
  assign binaryOp_40_io_enable_valid = bb_9_io_Out_2_valid; // @[bbgemm.scala 675:25]
  assign binaryOp_40_io_enable_bits_taskID = bb_9_io_Out_2_bits_taskID; // @[bbgemm.scala 675:25]
  assign binaryOp_40_io_enable_bits_control = bb_9_io_Out_2_bits_control; // @[bbgemm.scala 675:25]
  assign binaryOp_40_io_Out_0_ready = Loop_4_io_CarryDepenIn_0_ready; // @[bbgemm.scala 497:29]
  assign binaryOp_40_io_Out_1_ready = icmp_41_io_LeftIO_ready; // @[bbgemm.scala 843:21]
  assign binaryOp_40_io_LeftIO_valid = phi1_io_Out_1_valid; // @[bbgemm.scala 777:25]
  assign binaryOp_40_io_LeftIO_bits_taskID = phi1_io_Out_1_bits_taskID; // @[bbgemm.scala 777:25]
  assign binaryOp_40_io_LeftIO_bits_data = phi1_io_Out_1_bits_data; // @[bbgemm.scala 777:25]
  assign binaryOp_40_io_RightIO_valid = const15_io_Out_valid; // @[bbgemm.scala 773:26]
  assign binaryOp_40_io_RightIO_bits_taskID = const15_io_Out_bits_taskID; // @[bbgemm.scala 773:26]
  assign icmp_41_clock = clock;
  assign icmp_41_reset = reset;
  assign icmp_41_io_enable_valid = bb_9_io_Out_3_valid; // @[bbgemm.scala 678:21]
  assign icmp_41_io_enable_bits_taskID = bb_9_io_Out_3_bits_taskID; // @[bbgemm.scala 678:21]
  assign icmp_41_io_enable_bits_control = bb_9_io_Out_3_bits_control; // @[bbgemm.scala 678:21]
  assign icmp_41_io_Out_0_ready = br_42_io_CmpIO_ready; // @[bbgemm.scala 845:18]
  assign icmp_41_io_LeftIO_valid = binaryOp_40_io_Out_1_valid; // @[bbgemm.scala 843:21]
  assign icmp_41_io_LeftIO_bits_taskID = binaryOp_40_io_Out_1_bits_taskID; // @[bbgemm.scala 843:21]
  assign icmp_41_io_LeftIO_bits_data = binaryOp_40_io_Out_1_bits_data; // @[bbgemm.scala 843:21]
  assign icmp_41_io_RightIO_valid = const16_io_Out_valid; // @[bbgemm.scala 775:22]
  assign icmp_41_io_RightIO_bits_taskID = const16_io_Out_bits_taskID; // @[bbgemm.scala 775:22]
  assign br_42_clock = clock;
  assign br_42_reset = reset;
  assign br_42_io_enable_valid = bb_9_io_Out_4_valid; // @[bbgemm.scala 681:19]
  assign br_42_io_enable_bits_taskID = bb_9_io_Out_4_bits_taskID; // @[bbgemm.scala 681:19]
  assign br_42_io_enable_bits_control = bb_9_io_Out_4_bits_control; // @[bbgemm.scala 681:19]
  assign br_42_io_CmpIO_valid = icmp_41_io_Out_0_valid; // @[bbgemm.scala 845:18]
  assign br_42_io_CmpIO_bits_taskID = icmp_41_io_Out_0_bits_taskID; // @[bbgemm.scala 845:18]
  assign br_42_io_CmpIO_bits_data = icmp_41_io_Out_0_bits_data; // @[bbgemm.scala 845:18]
  assign br_42_io_TrueOutput_0_ready = Loop_4_io_loopBack_0_ready; // @[bbgemm.scala 379:25]
  assign br_42_io_FalseOutput_0_ready = Loop_4_io_loopFinish_0_ready; // @[bbgemm.scala 381:27]
  assign ret_43_clock = clock;
  assign ret_43_reset = reset;
  assign ret_43_io_In_enable_valid = bb_10_io_Out_0_valid; // @[bbgemm.scala 684:23]
  assign ret_43_io_In_enable_bits_taskID = bb_10_io_Out_0_bits_taskID; // @[bbgemm.scala 684:23]
  assign ret_43_io_In_enable_bits_control = bb_10_io_Out_0_bits_control; // @[bbgemm.scala 684:23]
  assign ret_43_io_Out_ready = io_out_ready; // @[bbgemm.scala 855:10]
  assign const0_clock = clock;
  assign const0_reset = reset;
  assign const0_io_enable_valid = bb_1_io_Out_0_valid; // @[bbgemm.scala 524:20]
  assign const0_io_enable_bits_taskID = bb_1_io_Out_0_bits_taskID; // @[bbgemm.scala 524:20]
  assign const0_io_Out_ready = phi1_io_InData_0_ready; // @[bbgemm.scala 743:21]
  assign const1_clock = clock;
  assign const1_reset = reset;
  assign const1_io_enable_valid = bb_2_io_Out_0_valid; // @[bbgemm.scala 532:20]
  assign const1_io_enable_bits_taskID = bb_2_io_Out_0_bits_taskID; // @[bbgemm.scala 532:20]
  assign const1_io_Out_ready = phi3_io_InData_0_ready; // @[bbgemm.scala 745:21]
  assign const2_clock = clock;
  assign const2_reset = reset;
  assign const2_io_enable_valid = bb_3_io_Out_0_valid; // @[bbgemm.scala 540:20]
  assign const2_io_enable_bits_taskID = bb_3_io_Out_0_bits_taskID; // @[bbgemm.scala 540:20]
  assign const2_io_Out_ready = phi5_io_InData_0_ready; // @[bbgemm.scala 747:21]
  assign const3_clock = clock;
  assign const3_reset = reset;
  assign const3_io_enable_valid = bb_3_io_Out_1_valid; // @[bbgemm.scala 542:20]
  assign const3_io_Out_ready = binaryOp_6_io_RightIO_ready; // @[bbgemm.scala 749:25]
  assign const4_clock = clock;
  assign const4_reset = reset;
  assign const4_io_enable_valid = bb_4_io_Out_0_valid; // @[bbgemm.scala 553:20]
  assign const4_io_enable_bits_taskID = bb_4_io_Out_0_bits_taskID; // @[bbgemm.scala 553:20]
  assign const4_io_Out_ready = phi8_io_InData_0_ready; // @[bbgemm.scala 751:21]
  assign const5_clock = clock;
  assign const5_reset = reset;
  assign const5_io_enable_valid = bb_4_io_Out_1_valid; // @[bbgemm.scala 555:20]
  assign const5_io_Out_ready = binaryOp_10_io_RightIO_ready; // @[bbgemm.scala 753:26]
  assign const6_clock = clock;
  assign const6_reset = reset;
  assign const6_io_enable_valid = bb_5_io_Out_0_valid; // @[bbgemm.scala 581:20]
  assign const6_io_enable_bits_taskID = bb_5_io_Out_0_bits_taskID; // @[bbgemm.scala 581:20]
  assign const6_io_Out_ready = phi16_io_InData_0_ready; // @[bbgemm.scala 755:22]
  assign const7_clock = clock;
  assign const7_reset = reset;
  assign const7_io_enable_valid = bb_5_io_Out_1_valid; // @[bbgemm.scala 583:20]
  assign const7_io_enable_bits_taskID = bb_5_io_Out_1_bits_taskID; // @[bbgemm.scala 583:20]
  assign const7_io_Out_ready = binaryOp_28_io_RightIO_ready; // @[bbgemm.scala 757:26]
  assign const8_clock = clock;
  assign const8_reset = reset;
  assign const8_io_enable_valid = bb_5_io_Out_2_valid; // @[bbgemm.scala 585:20]
  assign const8_io_enable_bits_taskID = bb_5_io_Out_2_bits_taskID; // @[bbgemm.scala 585:20]
  assign const8_io_Out_ready = icmp_29_io_RightIO_ready; // @[bbgemm.scala 759:22]
  assign const9_clock = clock;
  assign const9_reset = reset;
  assign const9_io_enable_valid = bb_6_io_Out_0_valid; // @[bbgemm.scala 632:20]
  assign const9_io_enable_bits_taskID = bb_6_io_Out_0_bits_taskID; // @[bbgemm.scala 632:20]
  assign const9_io_Out_ready = binaryOp_31_io_RightIO_ready; // @[bbgemm.scala 761:26]
  assign const10_clock = clock;
  assign const10_reset = reset;
  assign const10_io_enable_valid = bb_6_io_Out_1_valid; // @[bbgemm.scala 634:21]
  assign const10_io_enable_bits_taskID = bb_6_io_Out_1_bits_taskID; // @[bbgemm.scala 634:21]
  assign const10_io_Out_ready = icmp_32_io_RightIO_ready; // @[bbgemm.scala 763:22]
  assign const11_clock = clock;
  assign const11_reset = reset;
  assign const11_io_enable_valid = bb_7_io_Out_0_valid; // @[bbgemm.scala 645:21]
  assign const11_io_enable_bits_taskID = bb_7_io_Out_0_bits_taskID; // @[bbgemm.scala 645:21]
  assign const11_io_Out_ready = binaryOp_34_io_RightIO_ready; // @[bbgemm.scala 765:26]
  assign const12_clock = clock;
  assign const12_reset = reset;
  assign const12_io_enable_valid = bb_7_io_Out_1_valid; // @[bbgemm.scala 647:21]
  assign const12_io_enable_bits_taskID = bb_7_io_Out_1_bits_taskID; // @[bbgemm.scala 647:21]
  assign const12_io_Out_ready = icmp_35_io_RightIO_ready; // @[bbgemm.scala 767:22]
  assign const13_clock = clock;
  assign const13_reset = reset;
  assign const13_io_enable_valid = bb_8_io_Out_0_valid; // @[bbgemm.scala 658:21]
  assign const13_io_enable_bits_taskID = bb_8_io_Out_0_bits_taskID; // @[bbgemm.scala 658:21]
  assign const13_io_Out_ready = binaryOp_37_io_RightIO_ready; // @[bbgemm.scala 769:26]
  assign const14_clock = clock;
  assign const14_reset = reset;
  assign const14_io_enable_valid = bb_8_io_Out_1_valid; // @[bbgemm.scala 660:21]
  assign const14_io_enable_bits_taskID = bb_8_io_Out_1_bits_taskID; // @[bbgemm.scala 660:21]
  assign const14_io_Out_ready = icmp_38_io_RightIO_ready; // @[bbgemm.scala 771:22]
  assign const15_clock = clock;
  assign const15_reset = reset;
  assign const15_io_enable_valid = bb_9_io_Out_0_valid; // @[bbgemm.scala 671:21]
  assign const15_io_enable_bits_taskID = bb_9_io_Out_0_bits_taskID; // @[bbgemm.scala 671:21]
  assign const15_io_Out_ready = binaryOp_40_io_RightIO_ready; // @[bbgemm.scala 773:26]
  assign const16_clock = clock;
  assign const16_reset = reset;
  assign const16_io_enable_valid = bb_9_io_Out_1_valid; // @[bbgemm.scala 673:21]
  assign const16_io_enable_bits_taskID = bb_9_io_Out_1_bits_taskID; // @[bbgemm.scala 673:21]
  assign const16_io_Out_ready = icmp_41_io_RightIO_ready; // @[bbgemm.scala 775:22]
endmodule
